`timescale 1ns / 1ps

module tb_nebula_traffic_pattern();
  
  localparam int CLK_PERIOD = 10; // 100 MHz clock
  localparam int MESH_WIDTH = 8;
  localparam int MESH_HEIGHT = 8;
  localparam int NUM_NODES = MESH_WIDTH * MESH_HEIGHT;
  
  logic clk = 0;
  logic rst_n = 0;
  
  // Clock generation
  always #(CLK_PERIOD/2) clk = ~clk;
  
  // DUT instantiation
  nebula_top #(
    .MESH_WIDTH(MESH_WIDTH),
    .MESH_HEIGHT(MESH_HEIGHT)
  ) dut (
    .clk(clk),
    .rst_n(rst_n),
    // Other signals...
  );
  
  initial begin
    $dumpfile("nebula_traffic_pattern.vcd");
    $dumpvars(0, tb_nebula_traffic_pattern);
    
    // Reset sequence
    rst_n = 0;
    #(CLK_PERIOD * 5);
    rst_n = 1;
    #(CLK_PERIOD * 2);
    
    // Traffic injection based on generated pattern
    // Inject packets at cycle 0\n    // Packet 0: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 1: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 2: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 3: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 4: 8 -> 3 (AXI_WRITE)\n    inject_packet(8, 3, 64, "AXI_WRITE");\n    // Packet 5: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 6: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Packet 7: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Packet 8: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 1\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 1\n    // Packet 9: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 10: 12 -> 3 (AXI_WRITE)\n    inject_packet(12, 3, 64, "AXI_WRITE");\n    // Wait until cycle 2\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 2\n    // Packet 11: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 12: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 13: 9 -> 7 (AXI_WRITE)\n    inject_packet(9, 7, 64, "AXI_WRITE");\n    // Packet 14: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 15: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 3\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 3\n    // Packet 16: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 17: 1 -> 8 (AXI_WRITE)\n    inject_packet(1, 8, 64, "AXI_WRITE");\n    // Packet 18: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 19: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 20: 15 -> 2 (AXI_WRITE)\n    inject_packet(15, 2, 64, "AXI_WRITE");\n    // Wait until cycle 4\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 4\n    // Packet 21: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 22: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 23: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 24: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Packet 25: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 5\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 5\n    // Packet 26: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 27: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 28: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 29: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 30: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 31: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 6\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 6\n    // Packet 32: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 33: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Packet 34: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Packet 35: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Packet 36: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 7\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 7\n    // Packet 37: 1 -> 4 (AXI_WRITE)\n    inject_packet(1, 4, 64, "AXI_WRITE");\n    // Packet 38: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 39: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 40: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 41: 9 -> 11 (AXI_READ)\n    inject_packet(9, 11, 64, "AXI_READ");\n    // Packet 42: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Packet 43: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 44: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 8\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 8\n    // Packet 45: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 46: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 47: 6 -> 8 (AXI_WRITE)\n    inject_packet(6, 8, 64, "AXI_WRITE");\n    // Packet 48: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 49: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 50: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Packet 51: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Packet 52: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Wait until cycle 9\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 9\n    // Packet 53: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 54: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 55: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 56: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 57: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Packet 58: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 10\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 10\n    // Packet 59: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 60: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 61: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 62: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 63: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 64: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 65: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 66: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 11\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 11\n    // Packet 67: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 68: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 69: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 70: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Packet 71: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 72: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 73: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 74: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 12\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 12\n    // Packet 75: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 76: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 77: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 13\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 13\n    // Packet 78: 3 -> 2 (AXI_READ)\n    inject_packet(3, 2, 64, "AXI_READ");\n    // Packet 79: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 80: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 81: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 82: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Wait until cycle 14\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 14\n    // Packet 83: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 84: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 85: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 86: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 87: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Packet 88: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 15\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 15\n    // Packet 89: 1 -> 15 (AXI_WRITE)\n    inject_packet(1, 15, 64, "AXI_WRITE");\n    // Packet 90: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 91: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Wait until cycle 16\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 16\n    // Packet 92: 3 -> 8 (AXI_READ)\n    inject_packet(3, 8, 64, "AXI_READ");\n    // Packet 93: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 94: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 95: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Packet 96: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Wait until cycle 17\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 17\n    // Packet 97: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 98: 7 -> 13 (AXI_WRITE)\n    inject_packet(7, 13, 64, "AXI_WRITE");\n    // Packet 99: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Wait until cycle 18\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 18\n    // Packet 100: 8 -> 3 (AXI_WRITE)\n    inject_packet(8, 3, 64, "AXI_WRITE");\n    // Packet 101: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Packet 102: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Packet 103: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 19\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 19\n    // Packet 104: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 105: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 106: 9 -> 15 (AXI_WRITE)\n    inject_packet(9, 15, 64, "AXI_WRITE");\n    // Packet 107: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 20\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 20\n    // Packet 108: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 109: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 21\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 21\n    // Packet 110: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 111: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 112: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 113: 7 -> 9 (AXI_READ)\n    inject_packet(7, 9, 64, "AXI_READ");\n    // Packet 114: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 22\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 22\n    // Packet 115: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 116: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 117: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 118: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Packet 119: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Packet 120: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 23\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 23\n    // Packet 121: 1 -> 10 (AXI_READ)\n    inject_packet(1, 10, 64, "AXI_READ");\n    // Packet 122: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 123: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 24\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 24\n    // Packet 124: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 125: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 126: 13 -> 4 (AXI_WRITE)\n    inject_packet(13, 4, 64, "AXI_WRITE");\n    // Wait until cycle 25\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 25\n    // Packet 127: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Packet 128: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Wait until cycle 26\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 26\n    // Packet 129: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 130: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 131: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 132: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 133: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 134: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 135: 11 -> 0 (AXI_READ)\n    inject_packet(11, 0, 64, "AXI_READ");\n    // Packet 136: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Packet 137: 15 -> 0 (AXI_WRITE)\n    inject_packet(15, 0, 64, "AXI_WRITE");\n    // Wait until cycle 27\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 27\n    // Packet 138: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 139: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 140: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Packet 141: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Wait until cycle 28\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 28\n    // Packet 142: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 143: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Packet 144: 9 -> 2 (AXI_READ)\n    inject_packet(9, 2, 64, "AXI_READ");\n    // Packet 145: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 146: 13 -> 4 (AXI_WRITE)\n    inject_packet(13, 4, 64, "AXI_WRITE");\n    // Wait until cycle 29\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 29\n    // Packet 147: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Wait until cycle 30\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 30\n    // Packet 148: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 149: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 150: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 31\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 31\n    // Packet 151: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 152: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 153: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Wait until cycle 32\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 32\n    // Packet 154: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 155: 7 -> 9 (AXI_READ)\n    inject_packet(7, 9, 64, "AXI_READ");\n    // Packet 156: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 157: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Packet 158: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 33\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 33\n    // Packet 159: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 160: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 161: 7 -> 9 (AXI_READ)\n    inject_packet(7, 9, 64, "AXI_READ");\n    // Packet 162: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Wait until cycle 34\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 34\n    // Packet 163: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 164: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 35\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 35\n    // Packet 165: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Wait until cycle 36\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 36\n    // Packet 166: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 167: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 37\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 37\n    // Packet 168: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 169: 9 -> 13 (AXI_READ)\n    inject_packet(9, 13, 64, "AXI_READ");\n    // Packet 170: 10 -> 5 (AXI_WRITE)\n    inject_packet(10, 5, 64, "AXI_WRITE");\n    // Packet 171: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 172: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Wait until cycle 38\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 38\n    // Packet 173: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 174: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 175: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 176: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 177: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 178: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 179: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Packet 180: 15 -> 13 (AXI_WRITE)\n    inject_packet(15, 13, 64, "AXI_WRITE");\n    // Wait until cycle 39\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 39\n    // Packet 181: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 182: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 183: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Wait until cycle 40\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 40\n    // Packet 184: 3 -> 5 (AXI_WRITE)\n    inject_packet(3, 5, 64, "AXI_WRITE");\n    // Packet 185: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 186: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 187: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 188: 14 -> 12 (AXI_READ)\n    inject_packet(14, 12, 64, "AXI_READ");\n    // Wait until cycle 41\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 41\n    // Packet 189: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 190: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Packet 191: 14 -> 15 (AXI_WRITE)\n    inject_packet(14, 15, 64, "AXI_WRITE");\n    // Wait until cycle 42\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 42\n    // Packet 192: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 193: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 194: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Wait until cycle 43\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 43\n    // Packet 195: 3 -> 12 (AXI_WRITE)\n    inject_packet(3, 12, 64, "AXI_WRITE");\n    // Packet 196: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 197: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 198: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Packet 199: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 200: 13 -> 5 (AXI_READ)\n    inject_packet(13, 5, 64, "AXI_READ");\n    // Wait until cycle 44\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 44\n    // Packet 201: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 202: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 203: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 204: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 205: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Packet 206: 12 -> 4 (AXI_READ)\n    inject_packet(12, 4, 64, "AXI_READ");\n    // Packet 207: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Wait until cycle 45\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 45\n    // Packet 208: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 209: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 210: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 211: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 212: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 213: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Packet 214: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 46\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 46\n    // Packet 215: 0 -> 12 (AXI_READ)\n    inject_packet(0, 12, 64, "AXI_READ");\n    // Packet 216: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 217: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Packet 218: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Packet 219: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Wait until cycle 47\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 47\n    // Packet 220: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 221: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Packet 222: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Wait until cycle 48\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 48\n    // Packet 223: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 224: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 225: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 226: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 227: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Wait until cycle 49\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 49\n    // Packet 228: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 229: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 230: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 231: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 232: 9 -> 13 (AXI_READ)\n    inject_packet(9, 13, 64, "AXI_READ");\n    // Packet 233: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Packet 234: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Packet 235: 15 -> 4 (AXI_READ)\n    inject_packet(15, 4, 64, "AXI_READ");\n    // Wait until cycle 50\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 50\n    // Packet 236: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 237: 5 -> 9 (AXI_READ)\n    inject_packet(5, 9, 64, "AXI_READ");\n    // Packet 238: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 239: 12 -> 5 (AXI_WRITE)\n    inject_packet(12, 5, 64, "AXI_WRITE");\n    // Wait until cycle 51\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 51\n    // Packet 240: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 241: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 242: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 243: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 244: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Packet 245: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Wait until cycle 52\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 52\n    // Packet 246: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 247: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 248: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Wait until cycle 53\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 53\n    // Packet 249: 6 -> 8 (AXI_WRITE)\n    inject_packet(6, 8, 64, "AXI_WRITE");\n    // Packet 250: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 251: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Wait until cycle 54\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 54\n    // Packet 252: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 253: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 254: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 255: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Wait until cycle 55\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 55\n    // Packet 256: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 257: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 258: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 259: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Wait until cycle 56\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 56\n    // Packet 260: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 261: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 262: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Wait until cycle 57\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 57\n    // Packet 263: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 264: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 265: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Wait until cycle 58\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 58\n    // Packet 266: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 267: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 268: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 269: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Packet 270: 12 -> 13 (AXI_READ)\n    inject_packet(12, 13, 64, "AXI_READ");\n    // Packet 271: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 272: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 59\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 59\n    // Packet 273: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 274: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 275: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 276: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Packet 277: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 60\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 60\n    // Packet 278: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 279: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 280: 6 -> 7 (AXI_WRITE)\n    inject_packet(6, 7, 64, "AXI_WRITE");\n    // Packet 281: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 282: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 283: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Packet 284: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 285: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Wait until cycle 61\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 61\n    // Packet 286: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 287: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 288: 5 -> 0 (AXI_WRITE)\n    inject_packet(5, 0, 64, "AXI_WRITE");\n    // Packet 289: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Packet 290: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 62\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 62\n    // Packet 291: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 292: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 293: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 294: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Wait until cycle 63\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 63\n    // Packet 295: 1 -> 6 (AXI_WRITE)\n    inject_packet(1, 6, 64, "AXI_WRITE");\n    // Packet 296: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 64\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 64\n    // Packet 297: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 298: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Packet 299: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Wait until cycle 65\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 65\n    // Packet 300: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 301: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 302: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 66\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 66\n    // Packet 303: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 304: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 305: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 306: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Wait until cycle 67\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 67\n    // Packet 307: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 308: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 309: 7 -> 8 (AXI_READ)\n    inject_packet(7, 8, 64, "AXI_READ");\n    // Packet 310: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Packet 311: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Wait until cycle 68\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 68\n    // Packet 312: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 313: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 314: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 69\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 69\n    // Packet 315: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 316: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 317: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 318: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 319: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Wait until cycle 70\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 70\n    // Packet 320: 2 -> 5 (AXI_WRITE)\n    inject_packet(2, 5, 64, "AXI_WRITE");\n    // Packet 321: 3 -> 13 (AXI_WRITE)\n    inject_packet(3, 13, 64, "AXI_WRITE");\n    // Packet 322: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 323: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Packet 324: 8 -> 14 (AXI_WRITE)\n    inject_packet(8, 14, 64, "AXI_WRITE");\n    // Packet 325: 12 -> 5 (AXI_READ)\n    inject_packet(12, 5, 64, "AXI_READ");\n    // Packet 326: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 71\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 71\n    // Packet 327: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 328: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 329: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Packet 330: 15 -> 5 (AXI_READ)\n    inject_packet(15, 5, 64, "AXI_READ");\n    // Wait until cycle 72\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 72\n    // Packet 331: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 332: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 333: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 334: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 335: 12 -> 9 (AXI_READ)\n    inject_packet(12, 9, 64, "AXI_READ");\n    // Packet 336: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Wait until cycle 73\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 73\n    // Packet 337: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 338: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 339: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 340: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Wait until cycle 74\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 74\n    // Packet 341: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 342: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 343: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Packet 344: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 75\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 75\n    // Packet 345: 0 -> 12 (AXI_READ)\n    inject_packet(0, 12, 64, "AXI_READ");\n    // Packet 346: 1 -> 8 (AXI_WRITE)\n    inject_packet(1, 8, 64, "AXI_WRITE");\n    // Packet 347: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 348: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Wait until cycle 76\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 76\n    // Packet 349: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 350: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Wait until cycle 77\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 77\n    // Packet 351: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 352: 6 -> 0 (AXI_WRITE)\n    inject_packet(6, 0, 64, "AXI_WRITE");\n    // Packet 353: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 354: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 355: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Packet 356: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 78\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 78\n    // Packet 357: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 358: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 359: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 360: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 361: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 362: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 363: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 79\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 79\n    // Packet 364: 0 -> 14 (AXI_WRITE)\n    inject_packet(0, 14, 64, "AXI_WRITE");\n    // Packet 365: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 366: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 367: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 368: 12 -> 13 (AXI_READ)\n    inject_packet(12, 13, 64, "AXI_READ");\n    // Wait until cycle 80\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 80\n    // Packet 369: 1 -> 6 (AXI_WRITE)\n    inject_packet(1, 6, 64, "AXI_WRITE");\n    // Packet 370: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 371: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 372: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 373: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 374: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 375: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 81\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 81\n    // Packet 376: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 377: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 378: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 379: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Wait until cycle 82\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 82\n    // Packet 380: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 381: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 382: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 383: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 384: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 385: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 83\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 83\n    // Packet 386: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 387: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 388: 10 -> 2 (AXI_READ)\n    inject_packet(10, 2, 64, "AXI_READ");\n    // Wait until cycle 84\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 84\n    // Packet 389: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 390: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 85\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 85\n    // Packet 391: 2 -> 8 (AXI_WRITE)\n    inject_packet(2, 8, 64, "AXI_WRITE");\n    // Packet 392: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 393: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 394: 8 -> 1 (AXI_READ)\n    inject_packet(8, 1, 64, "AXI_READ");\n    // Packet 395: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 86\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 86\n    // Packet 396: 2 -> 5 (AXI_READ)\n    inject_packet(2, 5, 64, "AXI_READ");\n    // Packet 397: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 398: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Wait until cycle 87\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 87\n    // Packet 399: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Wait until cycle 88\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 88\n    // Packet 400: 1 -> 4 (AXI_WRITE)\n    inject_packet(1, 4, 64, "AXI_WRITE");\n    // Packet 401: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 402: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 403: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 404: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 405: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 406: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 89\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 89\n    // Packet 407: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 408: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 409: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Packet 410: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 90\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 90\n    // Packet 411: 1 -> 9 (AXI_WRITE)\n    inject_packet(1, 9, 64, "AXI_WRITE");\n    // Packet 412: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 413: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 414: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 415: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 416: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Packet 417: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 91\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 91\n    // Packet 418: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 419: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 420: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 421: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 422: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Packet 423: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 92\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 92\n    // Packet 424: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 425: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 426: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 427: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 428: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Wait until cycle 93\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 93\n    // Packet 429: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 430: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 431: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 432: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 433: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Packet 434: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Packet 435: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Wait until cycle 94\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 94\n    // Packet 436: 1 -> 3 (AXI_READ)\n    inject_packet(1, 3, 64, "AXI_READ");\n    // Packet 437: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Packet 438: 11 -> 6 (AXI_READ)\n    inject_packet(11, 6, 64, "AXI_READ");\n    // Wait until cycle 95\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 95\n    // Packet 439: 2 -> 5 (AXI_WRITE)\n    inject_packet(2, 5, 64, "AXI_WRITE");\n    // Packet 440: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 441: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Wait until cycle 96\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 96\n    // Packet 442: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 443: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 444: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 445: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Wait until cycle 97\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 97\n    // Packet 446: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 447: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 448: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 449: 6 -> 4 (AXI_WRITE)\n    inject_packet(6, 4, 64, "AXI_WRITE");\n    // Packet 450: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 451: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 98\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 98\n    // Packet 452: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 453: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 454: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Packet 455: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 99\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 99\n    // Packet 456: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 457: 8 -> 12 (AXI_READ)\n    inject_packet(8, 12, 64, "AXI_READ");\n    // Packet 458: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Wait until cycle 100\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 100\n    // Packet 459: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 460: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 461: 8 -> 3 (AXI_WRITE)\n    inject_packet(8, 3, 64, "AXI_WRITE");\n    // Packet 462: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Wait until cycle 101\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 101\n    // Packet 463: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 464: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 465: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 466: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Wait until cycle 102\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 102\n    // Packet 467: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 468: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 469: 8 -> 12 (AXI_READ)\n    inject_packet(8, 12, 64, "AXI_READ");\n    // Wait until cycle 103\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 103\n    // Packet 470: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 471: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 472: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 473: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Wait until cycle 104\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 104\n    // Packet 474: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 475: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 476: 10 -> 1 (AXI_READ)\n    inject_packet(10, 1, 64, "AXI_READ");\n    // Packet 477: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 105\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 105\n    // Packet 478: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 479: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 480: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Wait until cycle 106\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 106\n    // Packet 481: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 482: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 483: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 484: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 485: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 107\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 107\n    // Packet 486: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 487: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Wait until cycle 108\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 108\n    // Packet 488: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 489: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 490: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 491: 10 -> 14 (AXI_READ)\n    inject_packet(10, 14, 64, "AXI_READ");\n    // Packet 492: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Wait until cycle 109\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 109\n    // Packet 493: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 494: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 495: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Wait until cycle 110\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 110\n    // Packet 496: 5 -> 9 (AXI_READ)\n    inject_packet(5, 9, 64, "AXI_READ");\n    // Packet 497: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 498: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 499: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Wait until cycle 111\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 111\n    // Packet 500: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 501: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 502: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 503: 10 -> 1 (AXI_READ)\n    inject_packet(10, 1, 64, "AXI_READ");\n    // Packet 504: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 505: 15 -> 5 (AXI_READ)\n    inject_packet(15, 5, 64, "AXI_READ");\n    // Wait until cycle 112\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 112\n    // Packet 506: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 507: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 508: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 509: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 510: 12 -> 5 (AXI_READ)\n    inject_packet(12, 5, 64, "AXI_READ");\n    // Packet 511: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Wait until cycle 113\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 113\n    // Packet 512: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 513: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Packet 514: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Wait until cycle 114\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 114\n    // Packet 515: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 516: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 517: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 518: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Packet 519: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 115\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 115\n    // Packet 520: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 521: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 522: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 523: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Wait until cycle 116\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 116\n    // Packet 524: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 525: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 526: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 527: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 528: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 529: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Wait until cycle 117\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 117\n    // Packet 530: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 531: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 532: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 533: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 534: 7 -> 14 (AXI_READ)\n    inject_packet(7, 14, 64, "AXI_READ");\n    // Packet 535: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 536: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Wait until cycle 118\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 118\n    // Packet 537: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 538: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 539: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 540: 6 -> 8 (AXI_WRITE)\n    inject_packet(6, 8, 64, "AXI_WRITE");\n    // Packet 541: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 542: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 543: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Wait until cycle 119\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 119\n    // Packet 544: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 545: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 546: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 547: 12 -> 3 (AXI_WRITE)\n    inject_packet(12, 3, 64, "AXI_WRITE");\n    // Packet 548: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Packet 549: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 120\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 120\n    // Packet 550: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 551: 9 -> 11 (AXI_READ)\n    inject_packet(9, 11, 64, "AXI_READ");\n    // Packet 552: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Wait until cycle 121\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 121\n    // Packet 553: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 554: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 555: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 556: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 557: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Packet 558: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Packet 559: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 122\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 122\n    // Packet 560: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 561: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 562: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 563: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 564: 8 -> 14 (AXI_WRITE)\n    inject_packet(8, 14, 64, "AXI_WRITE");\n    // Packet 565: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Packet 566: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 123\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 123\n    // Packet 567: 1 -> 15 (AXI_WRITE)\n    inject_packet(1, 15, 64, "AXI_WRITE");\n    // Packet 568: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 569: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 570: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 571: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 572: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 573: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 574: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 124\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 124\n    // Packet 575: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 576: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 577: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Packet 578: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Wait until cycle 125\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 125\n    // Packet 579: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 580: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 581: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 582: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 126\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 126\n    // Packet 583: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 584: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 585: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 586: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 587: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 588: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Wait until cycle 127\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 127\n    // Packet 589: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 590: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 591: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 592: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 593: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 128\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 128\n    // Packet 594: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 595: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 596: 8 -> 12 (AXI_READ)\n    inject_packet(8, 12, 64, "AXI_READ");\n    // Packet 597: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Wait until cycle 129\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 129\n    // Packet 598: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 599: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 600: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 601: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Packet 602: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Packet 603: 15 -> 2 (AXI_WRITE)\n    inject_packet(15, 2, 64, "AXI_WRITE");\n    // Wait until cycle 130\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 130\n    // Packet 604: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 605: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Wait until cycle 131\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 131\n    // Packet 606: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 607: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 608: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 609: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 610: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 611: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Packet 612: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Packet 613: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Wait until cycle 132\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 132\n    // Packet 614: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 615: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 616: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 617: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 618: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 133\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 133\n    // Packet 619: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 620: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 621: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 622: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Packet 623: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 134\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 134\n    // Packet 624: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 625: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 626: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 627: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 135\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 135\n    // Packet 628: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 629: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 630: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Wait until cycle 136\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 136\n    // Packet 631: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 632: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 633: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Packet 634: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Packet 635: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Packet 636: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 137\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 137\n    // Packet 637: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 638: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 639: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 640: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 641: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 642: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 138\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 138\n    // Packet 643: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 644: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 645: 9 -> 2 (AXI_READ)\n    inject_packet(9, 2, 64, "AXI_READ");\n    // Packet 646: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Packet 647: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Wait until cycle 139\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 139\n    // Packet 648: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 649: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 650: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 651: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 652: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 653: 10 -> 8 (AXI_READ)\n    inject_packet(10, 8, 64, "AXI_READ");\n    // Wait until cycle 140\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 140\n    // Packet 654: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 655: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Packet 656: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 141\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 141\n    // Packet 657: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 658: 8 -> 3 (AXI_WRITE)\n    inject_packet(8, 3, 64, "AXI_WRITE");\n    // Packet 659: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 142\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 142\n    // Packet 660: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 661: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 662: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Packet 663: 15 -> 4 (AXI_READ)\n    inject_packet(15, 4, 64, "AXI_READ");\n    // Wait until cycle 143\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 143\n    // Packet 664: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 665: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 666: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 667: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Packet 668: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 144\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 144\n    // Packet 669: 1 -> 9 (AXI_WRITE)\n    inject_packet(1, 9, 64, "AXI_WRITE");\n    // Packet 670: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 671: 3 -> 5 (AXI_WRITE)\n    inject_packet(3, 5, 64, "AXI_WRITE");\n    // Packet 672: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 673: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Packet 674: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Packet 675: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 145\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 145\n    // Packet 676: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 677: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 678: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 679: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 680: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Wait until cycle 146\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 146\n    // Packet 681: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 682: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 683: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 147\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 147\n    // Packet 684: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 685: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 686: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Packet 687: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 148\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 148\n    // Packet 688: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 689: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 690: 7 -> 6 (AXI_WRITE)\n    inject_packet(7, 6, 64, "AXI_WRITE");\n    // Packet 691: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 692: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 693: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 149\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 149\n    // Packet 694: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 695: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Packet 696: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Wait until cycle 150\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 150\n    // Packet 697: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 698: 7 -> 14 (AXI_READ)\n    inject_packet(7, 14, 64, "AXI_READ");\n    // Packet 699: 8 -> 15 (AXI_READ)\n    inject_packet(8, 15, 64, "AXI_READ");\n    // Packet 700: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Packet 701: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 151\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 151\n    // Packet 702: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 703: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 704: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 705: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Wait until cycle 152\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 152\n    // Packet 706: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Packet 707: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Wait until cycle 153\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 153\n    // Packet 708: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 709: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 710: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Packet 711: 7 -> 14 (AXI_READ)\n    inject_packet(7, 14, 64, "AXI_READ");\n    // Packet 712: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Wait until cycle 154\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 154\n    // Packet 713: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 714: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 715: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 716: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Wait until cycle 155\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 155\n    // Packet 717: 0 -> 6 (AXI_WRITE)\n    inject_packet(0, 6, 64, "AXI_WRITE");\n    // Packet 718: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 719: 8 -> 3 (AXI_WRITE)\n    inject_packet(8, 3, 64, "AXI_WRITE");\n    // Packet 720: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 721: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 156\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 156\n    // Packet 722: 8 -> 1 (AXI_READ)\n    inject_packet(8, 1, 64, "AXI_READ");\n    // Packet 723: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 724: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Packet 725: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Packet 726: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 157\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 157\n    // Packet 727: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 728: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 729: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 730: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Packet 731: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Wait until cycle 158\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 158\n    // Packet 732: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 733: 9 -> 2 (AXI_READ)\n    inject_packet(9, 2, 64, "AXI_READ");\n    // Packet 734: 13 -> 9 (AXI_WRITE)\n    inject_packet(13, 9, 64, "AXI_WRITE");\n    // Packet 735: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Packet 736: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 159\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 159\n    // Packet 737: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Packet 738: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 739: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Wait until cycle 160\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 160\n    // Packet 740: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 741: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Wait until cycle 161\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 161\n    // Packet 742: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 743: 4 -> 11 (AXI_READ)\n    inject_packet(4, 11, 64, "AXI_READ");\n    // Packet 744: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 745: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 746: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Wait until cycle 162\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 162\n    // Packet 747: 2 -> 8 (AXI_WRITE)\n    inject_packet(2, 8, 64, "AXI_WRITE");\n    // Packet 748: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 749: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 750: 6 -> 4 (AXI_WRITE)\n    inject_packet(6, 4, 64, "AXI_WRITE");\n    // Packet 751: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Wait until cycle 163\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 163\n    // Packet 752: 1 -> 15 (AXI_READ)\n    inject_packet(1, 15, 64, "AXI_READ");\n    // Packet 753: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 754: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Packet 755: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Packet 756: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 757: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Packet 758: 12 -> 14 (AXI_READ)\n    inject_packet(12, 14, 64, "AXI_READ");\n    // Packet 759: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 164\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 164\n    // Packet 760: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Packet 761: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 762: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Packet 763: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 165\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 165\n    // Packet 764: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 765: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 166\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 166\n    // Packet 766: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 767: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 768: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Packet 769: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Wait until cycle 167\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 167\n    // Packet 770: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 771: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 772: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Wait until cycle 168\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 168\n    // Packet 773: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 774: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 775: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 776: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 777: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 778: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Packet 779: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 169\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 169\n    // Packet 780: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 781: 6 -> 4 (AXI_WRITE)\n    inject_packet(6, 4, 64, "AXI_WRITE");\n    // Packet 782: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 783: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 784: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 170\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 170\n    // Packet 785: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 786: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 787: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 788: 9 -> 0 (AXI_READ)\n    inject_packet(9, 0, 64, "AXI_READ");\n    // Packet 789: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 790: 13 -> 2 (AXI_WRITE)\n    inject_packet(13, 2, 64, "AXI_WRITE");\n    // Wait until cycle 171\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 171\n    // Packet 791: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 792: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 793: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Packet 794: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 172\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 172\n    // Packet 795: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 796: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 797: 8 -> 15 (AXI_READ)\n    inject_packet(8, 15, 64, "AXI_READ");\n    // Packet 798: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Packet 799: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 173\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 173\n    // Packet 800: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 801: 3 -> 13 (AXI_WRITE)\n    inject_packet(3, 13, 64, "AXI_WRITE");\n    // Packet 802: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 803: 12 -> 14 (AXI_READ)\n    inject_packet(12, 14, 64, "AXI_READ");\n    // Packet 804: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Packet 805: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 174\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 174\n    // Packet 806: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 807: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 808: 6 -> 9 (AXI_WRITE)\n    inject_packet(6, 9, 64, "AXI_WRITE");\n    // Packet 809: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 810: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 811: 13 -> 4 (AXI_WRITE)\n    inject_packet(13, 4, 64, "AXI_WRITE");\n    // Wait until cycle 175\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 175\n    // Packet 812: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 813: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 814: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 815: 14 -> 4 (AXI_READ)\n    inject_packet(14, 4, 64, "AXI_READ");\n    // Wait until cycle 176\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 176\n    // Packet 816: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 817: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Packet 818: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Wait until cycle 177\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 177\n    // Packet 819: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 820: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 821: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Wait until cycle 178\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 178\n    // Packet 822: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 823: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Wait until cycle 179\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 179\n    // Packet 824: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 825: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 826: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 827: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 828: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 829: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 830: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 180\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 180\n    // Packet 831: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 832: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 833: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 834: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Wait until cycle 181\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 181\n    // Packet 835: 4 -> 3 (AXI_READ)\n    inject_packet(4, 3, 64, "AXI_READ");\n    // Packet 836: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 837: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Packet 838: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 839: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 182\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 182\n    // Packet 840: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 841: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 842: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Wait until cycle 183\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 183\n    // Packet 843: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 844: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 845: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 846: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Wait until cycle 184\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 184\n    // Packet 847: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 848: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 849: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 850: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Wait until cycle 185\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 185\n    // Packet 851: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Wait until cycle 186\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 186\n    // Packet 852: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 853: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 854: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 855: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 856: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 857: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 858: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 859: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Packet 860: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Packet 861: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 187\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 187\n    // Packet 862: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 863: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Wait until cycle 188\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 188\n    // Packet 864: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 865: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 866: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 867: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 868: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 189\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 189\n    // Packet 869: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 870: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 871: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 872: 12 -> 4 (AXI_READ)\n    inject_packet(12, 4, 64, "AXI_READ");\n    // Packet 873: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 190\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 190\n    // Packet 874: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 875: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 876: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 877: 3 -> 12 (AXI_WRITE)\n    inject_packet(3, 12, 64, "AXI_WRITE");\n    // Packet 878: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Wait until cycle 191\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 191\n    // Packet 879: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 880: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 881: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 882: 5 -> 13 (AXI_READ)\n    inject_packet(5, 13, 64, "AXI_READ");\n    // Packet 883: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Wait until cycle 192\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 192\n    // Packet 884: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 885: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 886: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 887: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 888: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 889: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Packet 890: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Packet 891: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Wait until cycle 193\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 193\n    // Packet 892: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 893: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 894: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Packet 895: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 194\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 194\n    // Packet 896: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 897: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 898: 8 -> 9 (AXI_READ)\n    inject_packet(8, 9, 64, "AXI_READ");\n    // Wait until cycle 195\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 195\n    // Packet 899: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 900: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 901: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 902: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 903: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 904: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Packet 905: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 196\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 196\n    // Packet 906: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 907: 5 -> 15 (AXI_READ)\n    inject_packet(5, 15, 64, "AXI_READ");\n    // Wait until cycle 197\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 197\n    // Packet 908: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 909: 4 -> 3 (AXI_READ)\n    inject_packet(4, 3, 64, "AXI_READ");\n    // Packet 910: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 911: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Wait until cycle 198\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 198\n    // Packet 912: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Wait until cycle 199\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 199\n    // Packet 913: 0 -> 9 (AXI_READ)\n    inject_packet(0, 9, 64, "AXI_READ");\n    // Packet 914: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 915: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Packet 916: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Wait until cycle 200\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 200\n    // Packet 917: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 918: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 919: 6 -> 4 (AXI_WRITE)\n    inject_packet(6, 4, 64, "AXI_WRITE");\n    // Packet 920: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 921: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Wait until cycle 201\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 201\n    // Packet 922: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 923: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 924: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 925: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 202\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 202\n    // Packet 926: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 927: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 928: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 929: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 930: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Packet 931: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 203\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 203\n    // Packet 932: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 933: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 934: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Packet 935: 13 -> 5 (AXI_READ)\n    inject_packet(13, 5, 64, "AXI_READ");\n    // Wait until cycle 204\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 204\n    // Packet 936: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 937: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 938: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Wait until cycle 205\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 205\n    // Packet 939: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 940: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 941: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 942: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 943: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 944: 11 -> 6 (AXI_READ)\n    inject_packet(11, 6, 64, "AXI_READ");\n    // Packet 945: 15 -> 3 (AXI_WRITE)\n    inject_packet(15, 3, 64, "AXI_WRITE");\n    // Wait until cycle 206\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 206\n    // Packet 946: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 947: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 948: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 949: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Packet 950: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 207\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 207\n    // Packet 951: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 952: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 953: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Wait until cycle 208\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 208\n    // Packet 954: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 955: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 956: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 209\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 209\n    // Packet 957: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 958: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 959: 5 -> 0 (AXI_WRITE)\n    inject_packet(5, 0, 64, "AXI_WRITE");\n    // Packet 960: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 961: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 962: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 963: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Wait until cycle 210\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 210\n    // Packet 964: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 965: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 966: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Wait until cycle 211\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 211\n    // Packet 967: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 968: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 969: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 970: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 971: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 972: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Wait until cycle 212\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 212\n    // Packet 973: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 974: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 975: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 976: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 977: 9 -> 1 (AXI_WRITE)\n    inject_packet(9, 1, 64, "AXI_WRITE");\n    // Packet 978: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 979: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 213\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 213\n    // Packet 980: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 981: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 982: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 983: 10 -> 2 (AXI_READ)\n    inject_packet(10, 2, 64, "AXI_READ");\n    // Packet 984: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 985: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 986: 14 -> 15 (AXI_WRITE)\n    inject_packet(14, 15, 64, "AXI_WRITE");\n    // Packet 987: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 214\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 214\n    // Packet 988: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 989: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Packet 990: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 991: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Packet 992: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 993: 14 -> 4 (AXI_READ)\n    inject_packet(14, 4, 64, "AXI_READ");\n    // Wait until cycle 215\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 215\n    // Packet 994: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 995: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 996: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 997: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 998: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Wait until cycle 216\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 216\n    // Packet 999: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 1000: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 1001: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 1002: 12 -> 0 (AXI_WRITE)\n    inject_packet(12, 0, 64, "AXI_WRITE");\n    // Packet 1003: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Wait until cycle 217\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 217\n    // Packet 1004: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 1005: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 1006: 10 -> 5 (AXI_WRITE)\n    inject_packet(10, 5, 64, "AXI_WRITE");\n    // Packet 1007: 15 -> 13 (AXI_WRITE)\n    inject_packet(15, 13, 64, "AXI_WRITE");\n    // Wait until cycle 218\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 218\n    // Packet 1008: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 1009: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 1010: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 1011: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Wait until cycle 219\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 219\n    // Packet 1012: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 1013: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 1014: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 1015: 15 -> 4 (AXI_READ)\n    inject_packet(15, 4, 64, "AXI_READ");\n    // Wait until cycle 220\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 220\n    // Packet 1016: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 1017: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 1018: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 1019: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 1020: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Wait until cycle 221\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 221\n    // Packet 1021: 1 -> 15 (AXI_READ)\n    inject_packet(1, 15, 64, "AXI_READ");\n    // Packet 1022: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 1023: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 1024: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 1025: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Packet 1026: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 1027: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Packet 1028: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Packet 1029: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Packet 1030: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 222\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 222\n    // Packet 1031: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 1032: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 1033: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 1034: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 1035: 14 -> 12 (AXI_READ)\n    inject_packet(14, 12, 64, "AXI_READ");\n    // Wait until cycle 223\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 223\n    // Packet 1036: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 1037: 3 -> 5 (AXI_WRITE)\n    inject_packet(3, 5, 64, "AXI_WRITE");\n    // Packet 1038: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 1039: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Wait until cycle 224\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 224\n    // Packet 1040: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 1041: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Wait until cycle 225\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 225\n    // Packet 1042: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 1043: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 1044: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 226\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 226\n    // Packet 1045: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 1046: 10 -> 2 (AXI_READ)\n    inject_packet(10, 2, 64, "AXI_READ");\n    // Packet 1047: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Packet 1048: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Packet 1049: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 227\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 227\n    // Packet 1050: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 1051: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 1052: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 1053: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Wait until cycle 228\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 228\n    // Packet 1054: 1 -> 3 (AXI_WRITE)\n    inject_packet(1, 3, 64, "AXI_WRITE");\n    // Packet 1055: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 1056: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 1057: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 1058: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 1059: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Wait until cycle 229\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 229\n    // Packet 1060: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 1061: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 1062: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 230\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 230\n    // Packet 1063: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 1064: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 1065: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 1066: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 1067: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 231\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 231\n    // Packet 1068: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 1069: 8 -> 12 (AXI_READ)\n    inject_packet(8, 12, 64, "AXI_READ");\n    // Packet 1070: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 1071: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Packet 1072: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Wait until cycle 232\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 232\n    // Packet 1073: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 1074: 9 -> 2 (AXI_READ)\n    inject_packet(9, 2, 64, "AXI_READ");\n    // Wait until cycle 233\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 233\n    // Packet 1075: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 1076: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 1077: 2 -> 8 (AXI_WRITE)\n    inject_packet(2, 8, 64, "AXI_WRITE");\n    // Packet 1078: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 1079: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 1080: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 1081: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 234\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 234\n    // Packet 1082: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 1083: 12 -> 5 (AXI_READ)\n    inject_packet(12, 5, 64, "AXI_READ");\n    // Packet 1084: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Packet 1085: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 235\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 235\n    // Packet 1086: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 1087: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 1088: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 1089: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Packet 1090: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 236\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 236\n    // Packet 1091: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 1092: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 1093: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 1094: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 1095: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 1096: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 1097: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 1098: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Wait until cycle 237\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 237\n    // Packet 1099: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 1100: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 1101: 4 -> 11 (AXI_READ)\n    inject_packet(4, 11, 64, "AXI_READ");\n    // Packet 1102: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Wait until cycle 238\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 238\n    // Packet 1103: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 1104: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 1105: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 1106: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Wait until cycle 239\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 239\n    // Packet 1107: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 1108: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 1109: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 1110: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 1111: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Wait until cycle 240\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 240\n    // Packet 1112: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 1113: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 1114: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 1115: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 1116: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Packet 1117: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 241\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 241\n    // Packet 1118: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 1119: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 1120: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 1121: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 1122: 11 -> 0 (AXI_READ)\n    inject_packet(11, 0, 64, "AXI_READ");\n    // Packet 1123: 13 -> 2 (AXI_WRITE)\n    inject_packet(13, 2, 64, "AXI_WRITE");\n    // Packet 1124: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Wait until cycle 242\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 242\n    // Packet 1125: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 1126: 3 -> 8 (AXI_READ)\n    inject_packet(3, 8, 64, "AXI_READ");\n    // Packet 1127: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 1128: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Packet 1129: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 1130: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 243\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 243\n    // Packet 1131: 0 -> 14 (AXI_WRITE)\n    inject_packet(0, 14, 64, "AXI_WRITE");\n    // Packet 1132: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 1133: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 1134: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 1135: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 1136: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 1137: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Packet 1138: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 244\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 244\n    // Packet 1139: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 1140: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 1141: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 1142: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 1143: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 1144: 11 -> 3 (AXI_WRITE)\n    inject_packet(11, 3, 64, "AXI_WRITE");\n    // Packet 1145: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 1146: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 245\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 245\n    // Packet 1147: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 1148: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 1149: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 1150: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 1151: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 1152: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 1153: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 246\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 246\n    // Packet 1154: 0 -> 14 (AXI_WRITE)\n    inject_packet(0, 14, 64, "AXI_WRITE");\n    // Packet 1155: 2 -> 8 (AXI_WRITE)\n    inject_packet(2, 8, 64, "AXI_WRITE");\n    // Packet 1156: 3 -> 12 (AXI_WRITE)\n    inject_packet(3, 12, 64, "AXI_WRITE");\n    // Packet 1157: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 1158: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 1159: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Wait until cycle 247\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 247\n    // Packet 1160: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 1161: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 1162: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 1163: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1164: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Wait until cycle 248\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 248\n    // Packet 1165: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Packet 1166: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 1167: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Wait until cycle 249\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 249\n    // Packet 1168: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 1169: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 1170: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Wait until cycle 250\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 250\n    // Packet 1171: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Wait until cycle 251\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 251\n    // Packet 1172: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 1173: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 1174: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1175: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 1176: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 1177: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 252\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 252\n    // Packet 1178: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Wait until cycle 253\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 253\n    // Packet 1179: 0 -> 6 (AXI_WRITE)\n    inject_packet(0, 6, 64, "AXI_WRITE");\n    // Packet 1180: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 1181: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 1182: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 1183: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 1184: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 1185: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 254\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 254\n    // Packet 1186: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 1187: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 1188: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Wait until cycle 255\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 255\n    // Packet 1189: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 1190: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 1191: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 1192: 9 -> 15 (AXI_WRITE)\n    inject_packet(9, 15, 64, "AXI_WRITE");\n    // Packet 1193: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Wait until cycle 256\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 256\n    // Packet 1194: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 1195: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 1196: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Packet 1197: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 257\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 257\n    // Packet 1198: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 1199: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Wait until cycle 258\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 258\n    // Packet 1200: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 1201: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 1202: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 1203: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 1204: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 1205: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Wait until cycle 259\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 259\n    // Packet 1206: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 1207: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 1208: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 1209: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Wait until cycle 260\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 260\n    // Packet 1210: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 1211: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 1212: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 1213: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Wait until cycle 261\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 261\n    // Packet 1214: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 1215: 14 -> 2 (AXI_READ)\n    inject_packet(14, 2, 64, "AXI_READ");\n    // Wait until cycle 262\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 262\n    // Packet 1216: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Packet 1217: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 1218: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Packet 1219: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 263\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 263\n    // Packet 1220: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 1221: 4 -> 1 (AXI_WRITE)\n    inject_packet(4, 1, 64, "AXI_WRITE");\n    // Packet 1222: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 1223: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 1224: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Packet 1225: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 1226: 14 -> 8 (AXI_READ)\n    inject_packet(14, 8, 64, "AXI_READ");\n    // Wait until cycle 264\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 264\n    // Packet 1227: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 1228: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 1229: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 1230: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Wait until cycle 265\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 265\n    // Packet 1231: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 1232: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 1233: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 266\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 266\n    // Packet 1234: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 1235: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 1236: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Wait until cycle 267\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 267\n    // Packet 1237: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 1238: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 1239: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Packet 1240: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 1241: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 268\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 268\n    // Packet 1242: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 1243: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 1244: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Wait until cycle 269\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 269\n    // Packet 1245: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 1246: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 1247: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 1248: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Wait until cycle 270\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 270\n    // Packet 1249: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 1250: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 1251: 9 -> 0 (AXI_READ)\n    inject_packet(9, 0, 64, "AXI_READ");\n    // Packet 1252: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Wait until cycle 271\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 271\n    // Packet 1253: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 1254: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 1255: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 1256: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 1257: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Wait until cycle 272\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 272\n    // Packet 1258: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Wait until cycle 273\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 273\n    // Packet 1259: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 1260: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 1261: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 1262: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 1263: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Packet 1264: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Wait until cycle 274\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 274\n    // Packet 1265: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 1266: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 1267: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 1268: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Packet 1269: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Wait until cycle 275\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 275\n    // Packet 1270: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 1271: 1 -> 10 (AXI_READ)\n    inject_packet(1, 10, 64, "AXI_READ");\n    // Packet 1272: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 1273: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 1274: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 1275: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 1276: 12 -> 14 (AXI_READ)\n    inject_packet(12, 14, 64, "AXI_READ");\n    // Packet 1277: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 276\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 276\n    // Packet 1278: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 1279: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 1280: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 1281: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Wait until cycle 277\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 277\n    // Packet 1282: 3 -> 7 (AXI_READ)\n    inject_packet(3, 7, 64, "AXI_READ");\n    // Packet 1283: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 1284: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Wait until cycle 278\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 278\n    // Packet 1285: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 1286: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 1287: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 279\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 279\n    // Packet 1288: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1289: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 1290: 12 -> 14 (AXI_READ)\n    inject_packet(12, 14, 64, "AXI_READ");\n    // Wait until cycle 280\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 280\n    // Packet 1291: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Wait until cycle 281\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 281\n    // Packet 1292: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 1293: 3 -> 2 (AXI_READ)\n    inject_packet(3, 2, 64, "AXI_READ");\n    // Packet 1294: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 282\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 282\n    // Packet 1295: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 1296: 1 -> 15 (AXI_WRITE)\n    inject_packet(1, 15, 64, "AXI_WRITE");\n    // Packet 1297: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 1298: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 1299: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 1300: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Packet 1301: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Wait until cycle 283\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 283\n    // Packet 1302: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 1303: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 1304: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Packet 1305: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 1306: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Wait until cycle 284\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 284\n    // Packet 1307: 1 -> 3 (AXI_WRITE)\n    inject_packet(1, 3, 64, "AXI_WRITE");\n    // Packet 1308: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 1309: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 1310: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 1311: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 285\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 285\n    // Packet 1312: 6 -> 9 (AXI_WRITE)\n    inject_packet(6, 9, 64, "AXI_WRITE");\n    // Packet 1313: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 1314: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 1315: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Wait until cycle 286\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 286\n    // Packet 1316: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 1317: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 1318: 8 -> 14 (AXI_WRITE)\n    inject_packet(8, 14, 64, "AXI_WRITE");\n    // Packet 1319: 9 -> 2 (AXI_READ)\n    inject_packet(9, 2, 64, "AXI_READ");\n    // Packet 1320: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 1321: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 1322: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 287\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 287\n    // Packet 1323: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 1324: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 1325: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 1326: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 1327: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Packet 1328: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Wait until cycle 288\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 288\n    // Packet 1329: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 1330: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 1331: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Packet 1332: 15 -> 1 (AXI_WRITE)\n    inject_packet(15, 1, 64, "AXI_WRITE");\n    // Wait until cycle 289\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 289\n    // Packet 1333: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 1334: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 1335: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 1336: 3 -> 13 (AXI_WRITE)\n    inject_packet(3, 13, 64, "AXI_WRITE");\n    // Packet 1337: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 1338: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 1339: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Wait until cycle 290\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 290\n    // Packet 1340: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 1341: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Packet 1342: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 291\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 291\n    // Packet 1343: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Wait until cycle 292\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 292\n    // Packet 1344: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 1345: 1 -> 3 (AXI_WRITE)\n    inject_packet(1, 3, 64, "AXI_WRITE");\n    // Packet 1346: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 1347: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Packet 1348: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Packet 1349: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Packet 1350: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 293\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 293\n    // Packet 1351: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Packet 1352: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 1353: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 294\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 294\n    // Packet 1354: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 1355: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 1356: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Packet 1357: 10 -> 7 (AXI_READ)\n    inject_packet(10, 7, 64, "AXI_READ");\n    // Packet 1358: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 1359: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 295\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 295\n    // Packet 1360: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 1361: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 296\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 296\n    // Packet 1362: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 1363: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Wait until cycle 297\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 297\n    // Packet 1364: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Packet 1365: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 1366: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 1367: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 1368: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 1369: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 298\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 298\n    // Packet 1370: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 1371: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 1372: 15 -> 0 (AXI_WRITE)\n    inject_packet(15, 0, 64, "AXI_WRITE");\n    // Wait until cycle 299\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 299\n    // Packet 1373: 7 -> 9 (AXI_READ)\n    inject_packet(7, 9, 64, "AXI_READ");\n    // Packet 1374: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 1375: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 1376: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 300\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 300\n    // Packet 1377: 1 -> 4 (AXI_WRITE)\n    inject_packet(1, 4, 64, "AXI_WRITE");\n    // Packet 1378: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 1379: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 1380: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 1381: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 301\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 301\n    // Packet 1382: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 1383: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Packet 1384: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 302\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 302\n    // Packet 1385: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Wait until cycle 303\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 303\n    // Packet 1386: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 1387: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 1388: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Packet 1389: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 304\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 304\n    // Packet 1390: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 1391: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 1392: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 1393: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 1394: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 305\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 305\n    // Packet 1395: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 1396: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 1397: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Wait until cycle 306\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 306\n    // Packet 1398: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 1399: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 1400: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 307\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 307\n    // Packet 1401: 0 -> 14 (AXI_WRITE)\n    inject_packet(0, 14, 64, "AXI_WRITE");\n    // Packet 1402: 1 -> 6 (AXI_WRITE)\n    inject_packet(1, 6, 64, "AXI_WRITE");\n    // Packet 1403: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 1404: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 1405: 9 -> 15 (AXI_WRITE)\n    inject_packet(9, 15, 64, "AXI_WRITE");\n    // Packet 1406: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 1407: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 1408: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 308\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 308\n    // Packet 1409: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 1410: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 1411: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 1412: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Wait until cycle 309\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 309\n    // Packet 1413: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 1414: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 1415: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Packet 1416: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 310\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 310\n    // Packet 1417: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 1418: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 1419: 6 -> 0 (AXI_WRITE)\n    inject_packet(6, 0, 64, "AXI_WRITE");\n    // Packet 1420: 8 -> 1 (AXI_READ)\n    inject_packet(8, 1, 64, "AXI_READ");\n    // Packet 1421: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 1422: 11 -> 6 (AXI_READ)\n    inject_packet(11, 6, 64, "AXI_READ");\n    // Packet 1423: 12 -> 5 (AXI_READ)\n    inject_packet(12, 5, 64, "AXI_READ");\n    // Packet 1424: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 311\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 311\n    // Packet 1425: 4 -> 3 (AXI_READ)\n    inject_packet(4, 3, 64, "AXI_READ");\n    // Packet 1426: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 1427: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 312\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 312\n    // Packet 1428: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 1429: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 1430: 4 -> 11 (AXI_READ)\n    inject_packet(4, 11, 64, "AXI_READ");\n    // Packet 1431: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 1432: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 1433: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Packet 1434: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 313\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 313\n    // Packet 1435: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 1436: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 1437: 6 -> 2 (AXI_WRITE)\n    inject_packet(6, 2, 64, "AXI_WRITE");\n    // Packet 1438: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 1439: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 314\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 314\n    // Packet 1440: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 1441: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 1442: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 315\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 315\n    // Packet 1443: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 1444: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 1445: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 1446: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 1447: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 1448: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Packet 1449: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Packet 1450: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 316\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 316\n    // Packet 1451: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 1452: 1 -> 3 (AXI_READ)\n    inject_packet(1, 3, 64, "AXI_READ");\n    // Packet 1453: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 1454: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 1455: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 1456: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 1457: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 317\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 317\n    // Packet 1458: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 1459: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 1460: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 1461: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Packet 1462: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 318\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 318\n    // Packet 1463: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 1464: 4 -> 1 (AXI_WRITE)\n    inject_packet(4, 1, 64, "AXI_WRITE");\n    // Packet 1465: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 1466: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 1467: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 319\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 319\n    // Packet 1468: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 1469: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 1470: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 1471: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Packet 1472: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 1473: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 1474: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Packet 1475: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 320\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 320\n    // Packet 1476: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 1477: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 1478: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Packet 1479: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 1480: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Wait until cycle 321\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 321\n    // Packet 1481: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 1482: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 1483: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 1484: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 322\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 322\n    // Packet 1485: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 1486: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 1487: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 323\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 323\n    // Packet 1488: 2 -> 5 (AXI_READ)\n    inject_packet(2, 5, 64, "AXI_READ");\n    // Packet 1489: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 1490: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 1491: 9 -> 11 (AXI_READ)\n    inject_packet(9, 11, 64, "AXI_READ");\n    // Packet 1492: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Packet 1493: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 324\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 324\n    // Packet 1494: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 1495: 7 -> 6 (AXI_WRITE)\n    inject_packet(7, 6, 64, "AXI_WRITE");\n    // Packet 1496: 15 -> 2 (AXI_WRITE)\n    inject_packet(15, 2, 64, "AXI_WRITE");\n    // Wait until cycle 325\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 325\n    // Packet 1497: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 1498: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 1499: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Wait until cycle 326\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 326\n    // Packet 1500: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 1501: 1 -> 15 (AXI_READ)\n    inject_packet(1, 15, 64, "AXI_READ");\n    // Packet 1502: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 1503: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Packet 1504: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 1505: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 1506: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Wait until cycle 327\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 327\n    // Packet 1507: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 1508: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 1509: 5 -> 9 (AXI_READ)\n    inject_packet(5, 9, 64, "AXI_READ");\n    // Packet 1510: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 1511: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 1512: 10 -> 5 (AXI_WRITE)\n    inject_packet(10, 5, 64, "AXI_WRITE");\n    // Packet 1513: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 328\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 328\n    // Packet 1514: 3 -> 5 (AXI_WRITE)\n    inject_packet(3, 5, 64, "AXI_WRITE");\n    // Packet 1515: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 1516: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 329\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 329\n    // Packet 1517: 7 -> 13 (AXI_WRITE)\n    inject_packet(7, 13, 64, "AXI_WRITE");\n    // Packet 1518: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 1519: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 1520: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 330\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 330\n    // Packet 1521: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 1522: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 1523: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 331\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 331\n    // Packet 1524: 4 -> 11 (AXI_READ)\n    inject_packet(4, 11, 64, "AXI_READ");\n    // Packet 1525: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 1526: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 1527: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 1528: 12 -> 5 (AXI_WRITE)\n    inject_packet(12, 5, 64, "AXI_WRITE");\n    // Packet 1529: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 332\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 332\n    // Packet 1530: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 1531: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 1532: 11 -> 0 (AXI_READ)\n    inject_packet(11, 0, 64, "AXI_READ");\n    // Packet 1533: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 333\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 333\n    // Packet 1534: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 1535: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 1536: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Wait until cycle 334\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 334\n    // Packet 1537: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 1538: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 1539: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 1540: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 1541: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Packet 1542: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 335\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 335\n    // Packet 1543: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 1544: 8 -> 9 (AXI_READ)\n    inject_packet(8, 9, 64, "AXI_READ");\n    // Packet 1545: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 1546: 15 -> 1 (AXI_WRITE)\n    inject_packet(15, 1, 64, "AXI_WRITE");\n    // Wait until cycle 336\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 336\n    // Packet 1547: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 1548: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 1549: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 1550: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 1551: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Packet 1552: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Wait until cycle 337\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 337\n    // Packet 1553: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 1554: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 1555: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 1556: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 1557: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 1558: 11 -> 3 (AXI_READ)\n    inject_packet(11, 3, 64, "AXI_READ");\n    // Packet 1559: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Packet 1560: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Packet 1561: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 338\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 338\n    // Packet 1562: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 1563: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 1564: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Wait until cycle 339\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 339\n    // Packet 1565: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 1566: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 1567: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Packet 1568: 15 -> 2 (AXI_WRITE)\n    inject_packet(15, 2, 64, "AXI_WRITE");\n    // Wait until cycle 340\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 340\n    // Packet 1569: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 1570: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 1571: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 1572: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Wait until cycle 341\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 341\n    // Packet 1573: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 1574: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 1575: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 1576: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Packet 1577: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 1578: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 1579: 14 -> 2 (AXI_READ)\n    inject_packet(14, 2, 64, "AXI_READ");\n    // Wait until cycle 342\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 342\n    // Packet 1580: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 1581: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 1582: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Packet 1583: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 1584: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 343\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 343\n    // Packet 1585: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 1586: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 1587: 5 -> 15 (AXI_READ)\n    inject_packet(5, 15, 64, "AXI_READ");\n    // Packet 1588: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Wait until cycle 344\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 344\n    // Packet 1589: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 1590: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 1591: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 1592: 12 -> 0 (AXI_WRITE)\n    inject_packet(12, 0, 64, "AXI_WRITE");\n    // Wait until cycle 345\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 345\n    // Packet 1593: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 1594: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 1595: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 1596: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 1597: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Wait until cycle 346\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 346\n    // Packet 1598: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 1599: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 1600: 6 -> 2 (AXI_WRITE)\n    inject_packet(6, 2, 64, "AXI_WRITE");\n    // Packet 1601: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 1602: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 1603: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 347\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 347\n    // Packet 1604: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 1605: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 1606: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 1607: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 1608: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 1609: 8 -> 3 (AXI_WRITE)\n    inject_packet(8, 3, 64, "AXI_WRITE");\n    // Packet 1610: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 1611: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 348\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 348\n    // Packet 1612: 2 -> 8 (AXI_WRITE)\n    inject_packet(2, 8, 64, "AXI_WRITE");\n    // Packet 1613: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 1614: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 1615: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Wait until cycle 349\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 349\n    // Packet 1616: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 1617: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 1618: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 1619: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 1620: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Wait until cycle 350\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 350\n    // Packet 1621: 6 -> 7 (AXI_WRITE)\n    inject_packet(6, 7, 64, "AXI_WRITE");\n    // Packet 1622: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 351\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 351\n    // Packet 1623: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 1624: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 1625: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Packet 1626: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 1627: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Wait until cycle 352\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 352\n    // Packet 1628: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 1629: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Packet 1630: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Wait until cycle 353\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 353\n    // Packet 1631: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 1632: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 1633: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 354\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 354\n    // Packet 1634: 2 -> 5 (AXI_READ)\n    inject_packet(2, 5, 64, "AXI_READ");\n    // Packet 1635: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 1636: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 1637: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Packet 1638: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Packet 1639: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 355\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 355\n    // Packet 1640: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 1641: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 1642: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 356\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 356\n    // Packet 1643: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 1644: 6 -> 2 (AXI_WRITE)\n    inject_packet(6, 2, 64, "AXI_WRITE");\n    // Packet 1645: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 1646: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 1647: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 1648: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 357\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 357\n    // Packet 1649: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 1650: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 1651: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Wait until cycle 358\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 358\n    // Packet 1652: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 1653: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1654: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 1655: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Packet 1656: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 1657: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 359\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 359\n    // Packet 1658: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Packet 1659: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 1660: 11 -> 9 (AXI_READ)\n    inject_packet(11, 9, 64, "AXI_READ");\n    // Packet 1661: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 1662: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 1663: 15 -> 4 (AXI_READ)\n    inject_packet(15, 4, 64, "AXI_READ");\n    // Wait until cycle 360\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 360\n    // Packet 1664: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 1665: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Wait until cycle 361\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 361\n    // Packet 1666: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 1667: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 1668: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 1669: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 1670: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 1671: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 1672: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Packet 1673: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 362\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 362\n    // Packet 1674: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 1675: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 1676: 10 -> 4 (AXI_READ)\n    inject_packet(10, 4, 64, "AXI_READ");\n    // Packet 1677: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 363\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 363\n    // Packet 1678: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 1679: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 1680: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 1681: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 1682: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 1683: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Packet 1684: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Packet 1685: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 364\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 364\n    // Packet 1686: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 1687: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 1688: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 1689: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 1690: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 1691: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 365\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 365\n    // Packet 1692: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Wait until cycle 366\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 366\n    // Packet 1693: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Packet 1694: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Wait until cycle 367\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 367\n    // Packet 1695: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 1696: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 1697: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 1698: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 1699: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 368\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 368\n    // Packet 1700: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 1701: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 1702: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 1703: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 1704: 7 -> 6 (AXI_WRITE)\n    inject_packet(7, 6, 64, "AXI_WRITE");\n    // Packet 1705: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 1706: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 1707: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 1708: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Packet 1709: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 1710: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Wait until cycle 369\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 369\n    // Packet 1711: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Packet 1712: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 1713: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Packet 1714: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Wait until cycle 370\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 370\n    // Packet 1715: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 1716: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 1717: 4 -> 1 (AXI_WRITE)\n    inject_packet(4, 1, 64, "AXI_WRITE");\n    // Packet 1718: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 1719: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 1720: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 1721: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Packet 1722: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Packet 1723: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Packet 1724: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 371\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 371\n    // Packet 1725: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 1726: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 1727: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 1728: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 1729: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 372\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 372\n    // Packet 1730: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 1731: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 1732: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 1733: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 1734: 12 -> 4 (AXI_READ)\n    inject_packet(12, 4, 64, "AXI_READ");\n    // Packet 1735: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 373\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 373\n    // Packet 1736: 1 -> 15 (AXI_READ)\n    inject_packet(1, 15, 64, "AXI_READ");\n    // Packet 1737: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 1738: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 1739: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Wait until cycle 374\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 374\n    // Packet 1740: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 1741: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 1742: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Wait until cycle 375\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 375\n    // Packet 1743: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 1744: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 1745: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 1746: 10 -> 14 (AXI_READ)\n    inject_packet(10, 14, 64, "AXI_READ");\n    // Packet 1747: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 1748: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Packet 1749: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 1750: 15 -> 2 (AXI_WRITE)\n    inject_packet(15, 2, 64, "AXI_WRITE");\n    // Wait until cycle 376\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 376\n    // Packet 1751: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 1752: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 1753: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 1754: 9 -> 0 (AXI_READ)\n    inject_packet(9, 0, 64, "AXI_READ");\n    // Packet 1755: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 1756: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 377\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 377\n    // Packet 1757: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 1758: 2 -> 5 (AXI_READ)\n    inject_packet(2, 5, 64, "AXI_READ");\n    // Packet 1759: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 1760: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 1761: 10 -> 14 (AXI_READ)\n    inject_packet(10, 14, 64, "AXI_READ");\n    // Packet 1762: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 1763: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 378\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 378\n    // Packet 1764: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 1765: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 1766: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 1767: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 1768: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 1769: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 379\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 379\n    // Packet 1770: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 1771: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 1772: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Packet 1773: 12 -> 4 (AXI_READ)\n    inject_packet(12, 4, 64, "AXI_READ");\n    // Packet 1774: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 380\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 380\n    // Packet 1775: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 1776: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 1777: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 1778: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 1779: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 1780: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Packet 1781: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Wait until cycle 381\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 381\n    // Packet 1782: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 1783: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 1784: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 1785: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 1786: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 1787: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Packet 1788: 15 -> 5 (AXI_READ)\n    inject_packet(15, 5, 64, "AXI_READ");\n    // Wait until cycle 382\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 382\n    // Packet 1789: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 1790: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 1791: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Wait until cycle 383\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 383\n    // Packet 1792: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 1793: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 1794: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 1795: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Wait until cycle 384\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 384\n    // Packet 1796: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 1797: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 1798: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 1799: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1800: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 1801: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 1802: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 1803: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 1804: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 385\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 385\n    // Packet 1805: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 1806: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 1807: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 1808: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 1809: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Wait until cycle 386\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 386\n    // Packet 1810: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Packet 1811: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 1812: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Packet 1813: 10 -> 1 (AXI_READ)\n    inject_packet(10, 1, 64, "AXI_READ");\n    // Packet 1814: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 1815: 12 -> 4 (AXI_READ)\n    inject_packet(12, 4, 64, "AXI_READ");\n    // Packet 1816: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Wait until cycle 387\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 387\n    // Packet 1817: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 1818: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 1819: 10 -> 5 (AXI_WRITE)\n    inject_packet(10, 5, 64, "AXI_WRITE");\n    // Wait until cycle 388\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 388\n    // Packet 1820: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 1821: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 1822: 9 -> 2 (AXI_READ)\n    inject_packet(9, 2, 64, "AXI_READ");\n    // Packet 1823: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 1824: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Packet 1825: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 389\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 389\n    // Packet 1826: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 1827: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 1828: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 1829: 9 -> 0 (AXI_READ)\n    inject_packet(9, 0, 64, "AXI_READ");\n    // Wait until cycle 390\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 390\n    // Packet 1830: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 1831: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 1832: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 1833: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 1834: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Wait until cycle 391\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 391\n    // Packet 1835: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 1836: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 1837: 7 -> 14 (AXI_READ)\n    inject_packet(7, 14, 64, "AXI_READ");\n    // Packet 1838: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 1839: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Wait until cycle 392\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 392\n    // Packet 1840: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 1841: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 1842: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Packet 1843: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Wait until cycle 393\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 393\n    // Packet 1844: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 1845: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 1846: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 1847: 9 -> 1 (AXI_WRITE)\n    inject_packet(9, 1, 64, "AXI_WRITE");\n    // Packet 1848: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 1849: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 394\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 394\n    // Packet 1850: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 1851: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 1852: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 395\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 395\n    // Packet 1853: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 1854: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Wait until cycle 396\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 396\n    // Packet 1855: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 1856: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 1857: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 1858: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Wait until cycle 397\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 397\n    // Packet 1859: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 1860: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 1861: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 398\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 398\n    // Packet 1862: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 1863: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 1864: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Packet 1865: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Wait until cycle 399\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 399\n    // Packet 1866: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 1867: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 1868: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Wait until cycle 400\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 400\n    // Packet 1869: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 1870: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 1871: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 1872: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 1873: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 1874: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Wait until cycle 401\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 401\n    // Packet 1875: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 1876: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1877: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 1878: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 1879: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 402\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 402\n    // Packet 1880: 0 -> 9 (AXI_READ)\n    inject_packet(0, 9, 64, "AXI_READ");\n    // Packet 1881: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 1882: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 1883: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 1884: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 1885: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Packet 1886: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Wait until cycle 403\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 403\n    // Packet 1887: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 1888: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Packet 1889: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 1890: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 404\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 404\n    // Packet 1891: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 1892: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 1893: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 1894: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 1895: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 1896: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Wait until cycle 405\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 405\n    // Packet 1897: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Packet 1898: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 1899: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 1900: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 1901: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 1902: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 406\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 406\n    // Packet 1903: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 1904: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 1905: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 1906: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 1907: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Packet 1908: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Wait until cycle 407\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 407\n    // Packet 1909: 2 -> 5 (AXI_READ)\n    inject_packet(2, 5, 64, "AXI_READ");\n    // Packet 1910: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 1911: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Packet 1912: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Packet 1913: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 408\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 408\n    // Packet 1914: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 1915: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 1916: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 1917: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 1918: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Wait until cycle 409\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 409\n    // Packet 1919: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 1920: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 1921: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1922: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Packet 1923: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Packet 1924: 12 -> 4 (AXI_READ)\n    inject_packet(12, 4, 64, "AXI_READ");\n    // Packet 1925: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Packet 1926: 14 -> 2 (AXI_READ)\n    inject_packet(14, 2, 64, "AXI_READ");\n    // Wait until cycle 410\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 410\n    // Packet 1927: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 1928: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 1929: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Wait until cycle 411\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 411\n    // Packet 1930: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 1931: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 1932: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Wait until cycle 412\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 412\n    // Packet 1933: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 1934: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 1935: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 1936: 10 -> 7 (AXI_READ)\n    inject_packet(10, 7, 64, "AXI_READ");\n    // Packet 1937: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 1938: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 413\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 413\n    // Packet 1939: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 1940: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 1941: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 1942: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 1943: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Wait until cycle 414\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 414\n    // Packet 1944: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 1945: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 1946: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 1947: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 1948: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Packet 1949: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 1950: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Packet 1951: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 415\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 415\n    // Packet 1952: 0 -> 6 (AXI_WRITE)\n    inject_packet(0, 6, 64, "AXI_WRITE");\n    // Packet 1953: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 1954: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 1955: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 1956: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 1957: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 416\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 416\n    // Packet 1958: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 1959: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 1960: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 1961: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 1962: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 417\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 417\n    // Packet 1963: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 1964: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 1965: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 1966: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Wait until cycle 418\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 418\n    // Packet 1967: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 1968: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 1969: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 1970: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 1971: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Packet 1972: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Packet 1973: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 419\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 419\n    // Packet 1974: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 1975: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 1976: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 1977: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 1978: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 1979: 12 -> 0 (AXI_WRITE)\n    inject_packet(12, 0, 64, "AXI_WRITE");\n    // Packet 1980: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 420\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 420\n    // Packet 1981: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 1982: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 1983: 5 -> 13 (AXI_READ)\n    inject_packet(5, 13, 64, "AXI_READ");\n    // Packet 1984: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 1985: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 1986: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Wait until cycle 421\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 421\n    // Packet 1987: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 1988: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 1989: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Packet 1990: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 422\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 422\n    // Packet 1991: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 1992: 6 -> 4 (AXI_WRITE)\n    inject_packet(6, 4, 64, "AXI_WRITE");\n    // Packet 1993: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 1994: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 423\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 423\n    // Packet 1995: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 1996: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 1997: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 1998: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 1999: 9 -> 1 (AXI_WRITE)\n    inject_packet(9, 1, 64, "AXI_WRITE");\n    // Wait until cycle 424\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 424\n    // Packet 2000: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 2001: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Packet 2002: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 2003: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Packet 2004: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 425\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 425\n    // Packet 2005: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 2006: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 2007: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 2008: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 2009: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 2010: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Wait until cycle 426\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 426\n    // Packet 2011: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 2012: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 2013: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 2014: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Packet 2015: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 427\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 427\n    // Packet 2016: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 2017: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 2018: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 2019: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Packet 2020: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Packet 2021: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 428\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 428\n    // Packet 2022: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 2023: 1 -> 8 (AXI_WRITE)\n    inject_packet(1, 8, 64, "AXI_WRITE");\n    // Packet 2024: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 2025: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 2026: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 2027: 13 -> 2 (AXI_WRITE)\n    inject_packet(13, 2, 64, "AXI_WRITE");\n    // Packet 2028: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Wait until cycle 429\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 429\n    // Packet 2029: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 2030: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 2031: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 2032: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 2033: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Packet 2034: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Wait until cycle 430\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 430\n    // Packet 2035: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 2036: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 2037: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 2038: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 2039: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Wait until cycle 431\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 431\n    // Packet 2040: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 2041: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 2042: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 2043: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 2044: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 432\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 432\n    // Packet 2045: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 2046: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 2047: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 2048: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Packet 2049: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 433\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 433\n    // Packet 2050: 0 -> 12 (AXI_READ)\n    inject_packet(0, 12, 64, "AXI_READ");\n    // Packet 2051: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 2052: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 2053: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Packet 2054: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 2055: 10 -> 8 (AXI_READ)\n    inject_packet(10, 8, 64, "AXI_READ");\n    // Packet 2056: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 434\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 434\n    // Packet 2057: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 2058: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 2059: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 2060: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Packet 2061: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Packet 2062: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Wait until cycle 435\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 435\n    // Packet 2063: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 2064: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 2065: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 2066: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 2067: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 2068: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Wait until cycle 436\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 436\n    // Packet 2069: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 2070: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 2071: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Wait until cycle 437\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 437\n    // Packet 2072: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 2073: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 2074: 7 -> 3 (AXI_WRITE)\n    inject_packet(7, 3, 64, "AXI_WRITE");\n    // Wait until cycle 438\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 438\n    // Packet 2075: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 2076: 4 -> 0 (AXI_WRITE)\n    inject_packet(4, 0, 64, "AXI_WRITE");\n    // Packet 2077: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 2078: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 2079: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Packet 2080: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Packet 2081: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 439\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 439\n    // Packet 2082: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 2083: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 2084: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 2085: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 2086: 8 -> 14 (AXI_WRITE)\n    inject_packet(8, 14, 64, "AXI_WRITE");\n    // Packet 2087: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 2088: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 2089: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Packet 2090: 13 -> 9 (AXI_WRITE)\n    inject_packet(13, 9, 64, "AXI_WRITE");\n    // Wait until cycle 440\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 440\n    // Packet 2091: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 2092: 1 -> 6 (AXI_WRITE)\n    inject_packet(1, 6, 64, "AXI_WRITE");\n    // Packet 2093: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 2094: 11 -> 9 (AXI_READ)\n    inject_packet(11, 9, 64, "AXI_READ");\n    // Wait until cycle 441\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 441\n    // Packet 2095: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 2096: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 2097: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 442\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 442\n    // Packet 2098: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 2099: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 2100: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Wait until cycle 443\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 443\n    // Packet 2101: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 2102: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 2103: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 2104: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 2105: 15 -> 1 (AXI_WRITE)\n    inject_packet(15, 1, 64, "AXI_WRITE");\n    // Wait until cycle 444\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 444\n    // Packet 2106: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 2107: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 2108: 3 -> 2 (AXI_READ)\n    inject_packet(3, 2, 64, "AXI_READ");\n    // Packet 2109: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 2110: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 2111: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 445\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 445\n    // Packet 2112: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Packet 2113: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 446\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 446\n    // Packet 2114: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 2115: 10 -> 2 (AXI_READ)\n    inject_packet(10, 2, 64, "AXI_READ");\n    // Packet 2116: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Wait until cycle 447\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 447\n    // Packet 2117: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 2118: 2 -> 5 (AXI_WRITE)\n    inject_packet(2, 5, 64, "AXI_WRITE");\n    // Packet 2119: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 2120: 10 -> 3 (AXI_READ)\n    inject_packet(10, 3, 64, "AXI_READ");\n    // Packet 2121: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 2122: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 448\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 448\n    // Packet 2123: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2124: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 2125: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Packet 2126: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 2127: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Packet 2128: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Wait until cycle 449\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 449\n    // Packet 2129: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 2130: 4 -> 1 (AXI_WRITE)\n    inject_packet(4, 1, 64, "AXI_WRITE");\n    // Packet 2131: 5 -> 9 (AXI_READ)\n    inject_packet(5, 9, 64, "AXI_READ");\n    // Packet 2132: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 2133: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 2134: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Packet 2135: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Wait until cycle 450\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 450\n    // Packet 2136: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 2137: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 2138: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 2139: 10 -> 4 (AXI_READ)\n    inject_packet(10, 4, 64, "AXI_READ");\n    // Wait until cycle 451\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 451\n    // Packet 2140: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 2141: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 2142: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 2143: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Wait until cycle 452\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 452\n    // Packet 2144: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 2145: 3 -> 13 (AXI_WRITE)\n    inject_packet(3, 13, 64, "AXI_WRITE");\n    // Packet 2146: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 2147: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 2148: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 453\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 453\n    // Packet 2149: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 2150: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 2151: 13 -> 2 (AXI_WRITE)\n    inject_packet(13, 2, 64, "AXI_WRITE");\n    // Packet 2152: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 454\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 454\n    // Packet 2153: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 2154: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 2155: 7 -> 4 (AXI_WRITE)\n    inject_packet(7, 4, 64, "AXI_WRITE");\n    // Packet 2156: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 2157: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Wait until cycle 455\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 455\n    // Packet 2158: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 2159: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 2160: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 2161: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 2162: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 2163: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 456\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 456\n    // Packet 2164: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 2165: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 2166: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 2167: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 2168: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 2169: 15 -> 2 (AXI_WRITE)\n    inject_packet(15, 2, 64, "AXI_WRITE");\n    // Wait until cycle 457\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 457\n    // Packet 2170: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 2171: 5 -> 4 (AXI_WRITE)\n    inject_packet(5, 4, 64, "AXI_WRITE");\n    // Packet 2172: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Packet 2173: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Wait until cycle 458\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 458\n    // Packet 2174: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 2175: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Packet 2176: 7 -> 8 (AXI_READ)\n    inject_packet(7, 8, 64, "AXI_READ");\n    // Packet 2177: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 2178: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Packet 2179: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 2180: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Packet 2181: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 459\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 459\n    // Packet 2182: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 2183: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 2184: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 2185: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 2186: 10 -> 1 (AXI_READ)\n    inject_packet(10, 1, 64, "AXI_READ");\n    // Packet 2187: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 2188: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 460\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 460\n    // Packet 2189: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 2190: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 2191: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 2192: 8 -> 9 (AXI_READ)\n    inject_packet(8, 9, 64, "AXI_READ");\n    // Packet 2193: 9 -> 2 (AXI_READ)\n    inject_packet(9, 2, 64, "AXI_READ");\n    // Packet 2194: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 2195: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Wait until cycle 461\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 461\n    // Packet 2196: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 2197: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 2198: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 2199: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 2200: 7 -> 9 (AXI_WRITE)\n    inject_packet(7, 9, 64, "AXI_WRITE");\n    // Packet 2201: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 462\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 462\n    // Packet 2202: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 2203: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 463\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 463\n    // Packet 2204: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 2205: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 2206: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 2207: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 2208: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Wait until cycle 464\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 464\n    // Packet 2209: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 2210: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 2211: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 465\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 465\n    // Packet 2212: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 2213: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 2214: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 2215: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Wait until cycle 466\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 466\n    // Packet 2216: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 2217: 3 -> 8 (AXI_READ)\n    inject_packet(3, 8, 64, "AXI_READ");\n    // Packet 2218: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 2219: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 2220: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 2221: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 2222: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 467\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 467\n    // Packet 2223: 0 -> 6 (AXI_WRITE)\n    inject_packet(0, 6, 64, "AXI_WRITE");\n    // Packet 2224: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 2225: 10 -> 4 (AXI_READ)\n    inject_packet(10, 4, 64, "AXI_READ");\n    // Packet 2226: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 468\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 468\n    // Packet 2227: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 2228: 1 -> 6 (AXI_WRITE)\n    inject_packet(1, 6, 64, "AXI_WRITE");\n    // Packet 2229: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 2230: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 2231: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Packet 2232: 14 -> 12 (AXI_READ)\n    inject_packet(14, 12, 64, "AXI_READ");\n    // Packet 2233: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 469\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 469\n    // Packet 2234: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 2235: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 2236: 9 -> 7 (AXI_WRITE)\n    inject_packet(9, 7, 64, "AXI_WRITE");\n    // Packet 2237: 12 -> 5 (AXI_WRITE)\n    inject_packet(12, 5, 64, "AXI_WRITE");\n    // Packet 2238: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Wait until cycle 470\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 470\n    // Packet 2239: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 2240: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Wait until cycle 471\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 471\n    // Packet 2241: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 2242: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 2243: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 2244: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 2245: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 472\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 472\n    // Packet 2246: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 2247: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 2248: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 2249: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 2250: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Packet 2251: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 473\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 473\n    // Packet 2252: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 2253: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 2254: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Packet 2255: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 474\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 474\n    // Packet 2256: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 2257: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 2258: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 2259: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 2260: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 2261: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Packet 2262: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 475\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 475\n    // Packet 2263: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 2264: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 2265: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 2266: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Packet 2267: 15 -> 13 (AXI_WRITE)\n    inject_packet(15, 13, 64, "AXI_WRITE");\n    // Wait until cycle 476\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 476\n    // Packet 2268: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2269: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 2270: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 2271: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 2272: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 2273: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 2274: 10 -> 1 (AXI_READ)\n    inject_packet(10, 1, 64, "AXI_READ");\n    // Packet 2275: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 2276: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 477\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 477\n    // Packet 2277: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 2278: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 2279: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 2280: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 2281: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Wait until cycle 478\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 478\n    // Packet 2282: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 2283: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 2284: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 2285: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 2286: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 2287: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 2288: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 2289: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 479\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 479\n    // Packet 2290: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2291: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Packet 2292: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 480\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 480\n    // Packet 2293: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 2294: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 2295: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 2296: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 481\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 481\n    // Packet 2297: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 2298: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 2299: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 2300: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 2301: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Wait until cycle 482\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 482\n    // Packet 2302: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 2303: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 2304: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 2305: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 2306: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 2307: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Wait until cycle 483\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 483\n    // Packet 2308: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 2309: 6 -> 10 (AXI_WRITE)\n    inject_packet(6, 10, 64, "AXI_WRITE");\n    // Packet 2310: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Packet 2311: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 2312: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 2313: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 2314: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 484\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 484\n    // Packet 2315: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 2316: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 2317: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 2318: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 485\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 485\n    // Packet 2319: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 2320: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 2321: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Wait until cycle 486\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 486\n    // Packet 2322: 1 -> 4 (AXI_WRITE)\n    inject_packet(1, 4, 64, "AXI_WRITE");\n    // Packet 2323: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 2324: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Packet 2325: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 2326: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 2327: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Wait until cycle 487\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 487\n    // Packet 2328: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 2329: 7 -> 4 (AXI_WRITE)\n    inject_packet(7, 4, 64, "AXI_WRITE");\n    // Packet 2330: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Packet 2331: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Wait until cycle 488\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 488\n    // Packet 2332: 15 -> 3 (AXI_WRITE)\n    inject_packet(15, 3, 64, "AXI_WRITE");\n    // Wait until cycle 489\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 489\n    // Packet 2333: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 2334: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 2335: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 2336: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 2337: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Packet 2338: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 490\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 490\n    // Packet 2339: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 2340: 3 -> 12 (AXI_WRITE)\n    inject_packet(3, 12, 64, "AXI_WRITE");\n    // Packet 2341: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 2342: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 2343: 8 -> 4 (AXI_READ)\n    inject_packet(8, 4, 64, "AXI_READ");\n    // Packet 2344: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 2345: 15 -> 1 (AXI_WRITE)\n    inject_packet(15, 1, 64, "AXI_WRITE");\n    // Wait until cycle 491\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 491\n    // Packet 2346: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 2347: 2 -> 8 (AXI_WRITE)\n    inject_packet(2, 8, 64, "AXI_WRITE");\n    // Packet 2348: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 2349: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Packet 2350: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 2351: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 2352: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 492\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 492\n    // Packet 2353: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 2354: 9 -> 1 (AXI_WRITE)\n    inject_packet(9, 1, 64, "AXI_WRITE");\n    // Packet 2355: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 2356: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 493\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 493\n    // Packet 2357: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 2358: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 2359: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 2360: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 2361: 14 -> 15 (AXI_WRITE)\n    inject_packet(14, 15, 64, "AXI_WRITE");\n    // Wait until cycle 494\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 494\n    // Packet 2362: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 2363: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 2364: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Packet 2365: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 495\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 495\n    // Packet 2366: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 2367: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 2368: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 2369: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Wait until cycle 496\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 496\n    // Packet 2370: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2371: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 2372: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 2373: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 2374: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Wait until cycle 497\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 497\n    // Packet 2375: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 2376: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 2377: 12 -> 5 (AXI_WRITE)\n    inject_packet(12, 5, 64, "AXI_WRITE");\n    // Packet 2378: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Packet 2379: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Packet 2380: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 498\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 498\n    // Packet 2381: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 2382: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 2383: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Wait until cycle 499\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 499\n    // Packet 2384: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 2385: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 2386: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Wait until cycle 500\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 500\n    // Packet 2387: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2388: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 2389: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 2390: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 2391: 11 -> 2 (AXI_READ)\n    inject_packet(11, 2, 64, "AXI_READ");\n    // Packet 2392: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Wait until cycle 501\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 501\n    // Packet 2393: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 2394: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Packet 2395: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 2396: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Wait until cycle 502\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 502\n    // Packet 2397: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 2398: 1 -> 3 (AXI_READ)\n    inject_packet(1, 3, 64, "AXI_READ");\n    // Packet 2399: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 2400: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 2401: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 503\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 503\n    // Packet 2402: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 2403: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 2404: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 2405: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 2406: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 2407: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Wait until cycle 504\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 504\n    // Packet 2408: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 2409: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 2410: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 2411: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Packet 2412: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 505\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 505\n    // Packet 2413: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 2414: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 2415: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 2416: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 2417: 12 -> 9 (AXI_READ)\n    inject_packet(12, 9, 64, "AXI_READ");\n    // Wait until cycle 506\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 506\n    // Packet 2418: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 2419: 3 -> 8 (AXI_READ)\n    inject_packet(3, 8, 64, "AXI_READ");\n    // Packet 2420: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 2421: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 2422: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 2423: 10 -> 4 (AXI_READ)\n    inject_packet(10, 4, 64, "AXI_READ");\n    // Wait until cycle 507\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 507\n    // Packet 2424: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 2425: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 2426: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 2427: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Packet 2428: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Wait until cycle 508\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 508\n    // Packet 2429: 0 -> 14 (AXI_WRITE)\n    inject_packet(0, 14, 64, "AXI_WRITE");\n    // Packet 2430: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 2431: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 2432: 7 -> 13 (AXI_WRITE)\n    inject_packet(7, 13, 64, "AXI_WRITE");\n    // Packet 2433: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 2434: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Packet 2435: 14 -> 8 (AXI_READ)\n    inject_packet(14, 8, 64, "AXI_READ");\n    // Packet 2436: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 509\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 509\n    // Packet 2437: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 2438: 1 -> 6 (AXI_WRITE)\n    inject_packet(1, 6, 64, "AXI_WRITE");\n    // Packet 2439: 7 -> 14 (AXI_READ)\n    inject_packet(7, 14, 64, "AXI_READ");\n    // Packet 2440: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 2441: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Packet 2442: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 510\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 510\n    // Packet 2443: 3 -> 2 (AXI_READ)\n    inject_packet(3, 2, 64, "AXI_READ");\n    // Packet 2444: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 2445: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Packet 2446: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 2447: 15 -> 4 (AXI_READ)\n    inject_packet(15, 4, 64, "AXI_READ");\n    // Wait until cycle 511\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 511\n    // Packet 2448: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 2449: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 2450: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 2451: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 2452: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 2453: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 2454: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 2455: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Packet 2456: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 512\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 512\n    // Packet 2457: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 2458: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 2459: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 2460: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 2461: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Wait until cycle 513\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 513\n    // Packet 2462: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 2463: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 514\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 514\n    // Packet 2464: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 2465: 4 -> 12 (AXI_WRITE)\n    inject_packet(4, 12, 64, "AXI_WRITE");\n    // Packet 2466: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 2467: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Wait until cycle 515\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 515\n    // Packet 2468: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Wait until cycle 516\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 516\n    // Packet 2469: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 2470: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 2471: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 2472: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 2473: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Wait until cycle 517\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 517\n    // Packet 2474: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 2475: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 2476: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 2477: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Wait until cycle 518\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 518\n    // Packet 2478: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 2479: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 2480: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Wait until cycle 519\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 519\n    // Packet 2481: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 2482: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 2483: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 2484: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 2485: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 2486: 11 -> 3 (AXI_READ)\n    inject_packet(11, 3, 64, "AXI_READ");\n    // Packet 2487: 12 -> 3 (AXI_WRITE)\n    inject_packet(12, 3, 64, "AXI_WRITE");\n    // Packet 2488: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Packet 2489: 15 -> 0 (AXI_WRITE)\n    inject_packet(15, 0, 64, "AXI_WRITE");\n    // Wait until cycle 520\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 520\n    // Packet 2490: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Wait until cycle 521\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 521\n    // Packet 2491: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 2492: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 2493: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Wait until cycle 522\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 522\n    // Packet 2494: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2495: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 2496: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 2497: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 2498: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Wait until cycle 523\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 523\n    // Packet 2499: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 2500: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 2501: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Wait until cycle 524\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 524\n    // Packet 2502: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 2503: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 2504: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 2505: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 2506: 13 -> 4 (AXI_WRITE)\n    inject_packet(13, 4, 64, "AXI_WRITE");\n    // Packet 2507: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Wait until cycle 525\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 525\n    // Packet 2508: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 2509: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 2510: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 2511: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 2512: 8 -> 9 (AXI_READ)\n    inject_packet(8, 9, 64, "AXI_READ");\n    // Packet 2513: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 2514: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 2515: 13 -> 9 (AXI_WRITE)\n    inject_packet(13, 9, 64, "AXI_WRITE");\n    // Packet 2516: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Packet 2517: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 526\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 526\n    // Packet 2518: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 2519: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 2520: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 2521: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Packet 2522: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Wait until cycle 527\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 527\n    // Packet 2523: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 2524: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 2525: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 2526: 14 -> 8 (AXI_READ)\n    inject_packet(14, 8, 64, "AXI_READ");\n    // Wait until cycle 528\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 528\n    // Packet 2527: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 2528: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Wait until cycle 529\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 529\n    // Packet 2529: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 2530: 4 -> 1 (AXI_WRITE)\n    inject_packet(4, 1, 64, "AXI_WRITE");\n    // Packet 2531: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 2532: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 2533: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Wait until cycle 530\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 530\n    // Packet 2534: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 2535: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 2536: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 2537: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 2538: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 2539: 10 -> 4 (AXI_READ)\n    inject_packet(10, 4, 64, "AXI_READ");\n    // Packet 2540: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 531\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 531\n    // Packet 2541: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 2542: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Packet 2543: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Wait until cycle 532\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 532\n    // Packet 2544: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 2545: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 2546: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 2547: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 2548: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 2549: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 2550: 6 -> 9 (AXI_WRITE)\n    inject_packet(6, 9, 64, "AXI_WRITE");\n    // Packet 2551: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Packet 2552: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 2553: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Wait until cycle 533\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 533\n    // Packet 2554: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 2555: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 2556: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 2557: 5 -> 13 (AXI_READ)\n    inject_packet(5, 13, 64, "AXI_READ");\n    // Packet 2558: 6 -> 10 (AXI_WRITE)\n    inject_packet(6, 10, 64, "AXI_WRITE");\n    // Packet 2559: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 2560: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 534\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 534\n    // Packet 2561: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 2562: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 2563: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 2564: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 2565: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 2566: 15 -> 1 (AXI_WRITE)\n    inject_packet(15, 1, 64, "AXI_WRITE");\n    // Wait until cycle 535\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 535\n    // Packet 2567: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 2568: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 2569: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 2570: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 2571: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Packet 2572: 14 -> 9 (AXI_WRITE)\n    inject_packet(14, 9, 64, "AXI_WRITE");\n    // Wait until cycle 536\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 536\n    // Packet 2573: 7 -> 9 (AXI_WRITE)\n    inject_packet(7, 9, 64, "AXI_WRITE");\n    // Packet 2574: 8 -> 4 (AXI_READ)\n    inject_packet(8, 4, 64, "AXI_READ");\n    // Packet 2575: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 2576: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 537\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 537\n    // Packet 2577: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 2578: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 2579: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Packet 2580: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Wait until cycle 539\n    repeat(2) @(posedge clk);\n    // Inject packets at cycle 539\n    // Packet 2581: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 2582: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 2583: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 2584: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 2585: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Wait until cycle 540\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 540\n    // Packet 2586: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 2587: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 2588: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 2589: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Packet 2590: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 2591: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 541\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 541\n    // Packet 2592: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 2593: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 2594: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 2595: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 2596: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 2597: 12 -> 0 (AXI_WRITE)\n    inject_packet(12, 0, 64, "AXI_WRITE");\n    // Packet 2598: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 542\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 542\n    // Packet 2599: 6 -> 2 (AXI_WRITE)\n    inject_packet(6, 2, 64, "AXI_WRITE");\n    // Packet 2600: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 2601: 14 -> 9 (AXI_WRITE)\n    inject_packet(14, 9, 64, "AXI_WRITE");\n    // Packet 2602: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 543\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 543\n    // Packet 2603: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 2604: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 2605: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 2606: 7 -> 6 (AXI_WRITE)\n    inject_packet(7, 6, 64, "AXI_WRITE");\n    // Packet 2607: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 2608: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Packet 2609: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Wait until cycle 544\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 544\n    // Packet 2610: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 2611: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 2612: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 545\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 545\n    // Packet 2613: 1 -> 3 (AXI_READ)\n    inject_packet(1, 3, 64, "AXI_READ");\n    // Packet 2614: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 2615: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 2616: 6 -> 0 (AXI_WRITE)\n    inject_packet(6, 0, 64, "AXI_WRITE");\n    // Packet 2617: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 2618: 14 -> 2 (AXI_READ)\n    inject_packet(14, 2, 64, "AXI_READ");\n    // Wait until cycle 546\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 546\n    // Packet 2619: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 2620: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 2621: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 2622: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Wait until cycle 547\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 547\n    // Packet 2623: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Packet 2624: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 2625: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 2626: 6 -> 7 (AXI_WRITE)\n    inject_packet(6, 7, 64, "AXI_WRITE");\n    // Packet 2627: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 2628: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 548\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 548\n    // Packet 2629: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 2630: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 2631: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Wait until cycle 549\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 549\n    // Packet 2632: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Wait until cycle 550\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 550\n    // Packet 2633: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 2634: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 2635: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 2636: 10 -> 2 (AXI_READ)\n    inject_packet(10, 2, 64, "AXI_READ");\n    // Packet 2637: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 2638: 12 -> 5 (AXI_READ)\n    inject_packet(12, 5, 64, "AXI_READ");\n    // Packet 2639: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Wait until cycle 551\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 551\n    // Packet 2640: 1 -> 8 (AXI_WRITE)\n    inject_packet(1, 8, 64, "AXI_WRITE");\n    // Packet 2641: 4 -> 11 (AXI_READ)\n    inject_packet(4, 11, 64, "AXI_READ");\n    // Packet 2642: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 2643: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 2644: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Wait until cycle 552\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 552\n    // Packet 2645: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 2646: 6 -> 8 (AXI_WRITE)\n    inject_packet(6, 8, 64, "AXI_WRITE");\n    // Packet 2647: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 2648: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Wait until cycle 553\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 553\n    // Packet 2649: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 2650: 13 -> 5 (AXI_READ)\n    inject_packet(13, 5, 64, "AXI_READ");\n    // Wait until cycle 554\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 554\n    // Packet 2651: 3 -> 7 (AXI_READ)\n    inject_packet(3, 7, 64, "AXI_READ");\n    // Packet 2652: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 2653: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 2654: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Wait until cycle 555\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 555\n    // Packet 2655: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 2656: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 2657: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 2658: 6 -> 7 (AXI_WRITE)\n    inject_packet(6, 7, 64, "AXI_WRITE");\n    // Packet 2659: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 2660: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 2661: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 2662: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 2663: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 556\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 556\n    // Packet 2664: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 2665: 1 -> 10 (AXI_READ)\n    inject_packet(1, 10, 64, "AXI_READ");\n    // Packet 2666: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 2667: 14 -> 4 (AXI_WRITE)\n    inject_packet(14, 4, 64, "AXI_WRITE");\n    // Wait until cycle 557\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 557\n    // Packet 2668: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 2669: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 2670: 7 -> 13 (AXI_WRITE)\n    inject_packet(7, 13, 64, "AXI_WRITE");\n    // Wait until cycle 558\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 558\n    // Packet 2671: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 2672: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Packet 2673: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 2674: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 2675: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 2676: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Wait until cycle 559\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 559\n    // Packet 2677: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 2678: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 2679: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 2680: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 2681: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Packet 2682: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 2683: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Wait until cycle 560\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 560\n    // Packet 2684: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 2685: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 2686: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 2687: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Wait until cycle 561\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 561\n    // Packet 2688: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 2689: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 2690: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 2691: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Wait until cycle 562\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 562\n    // Packet 2692: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 2693: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 2694: 11 -> 3 (AXI_WRITE)\n    inject_packet(11, 3, 64, "AXI_WRITE");\n    // Packet 2695: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Packet 2696: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 563\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 563\n    // Packet 2697: 1 -> 15 (AXI_READ)\n    inject_packet(1, 15, 64, "AXI_READ");\n    // Packet 2698: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 2699: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 2700: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 2701: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 2702: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Packet 2703: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Wait until cycle 564\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 564\n    // Packet 2704: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 2705: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 2706: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 2707: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Wait until cycle 565\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 565\n    // Packet 2708: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 2709: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 2710: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 566\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 566\n    // Packet 2711: 2 -> 5 (AXI_READ)\n    inject_packet(2, 5, 64, "AXI_READ");\n    // Packet 2712: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 2713: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 567\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 567\n    // Packet 2714: 10 -> 8 (AXI_READ)\n    inject_packet(10, 8, 64, "AXI_READ");\n    // Wait until cycle 568\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 568\n    // Packet 2715: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 2716: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 2717: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Wait until cycle 569\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 569\n    // Packet 2718: 4 -> 11 (AXI_READ)\n    inject_packet(4, 11, 64, "AXI_READ");\n    // Packet 2719: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 2720: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 2721: 10 -> 7 (AXI_READ)\n    inject_packet(10, 7, 64, "AXI_READ");\n    // Wait until cycle 570\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 570\n    // Packet 2722: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 2723: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Wait until cycle 571\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 571\n    // Packet 2724: 4 -> 5 (AXI_READ)\n    inject_packet(4, 5, 64, "AXI_READ");\n    // Packet 2725: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 2726: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 2727: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Wait until cycle 572\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 572\n    // Packet 2728: 1 -> 9 (AXI_WRITE)\n    inject_packet(1, 9, 64, "AXI_WRITE");\n    // Packet 2729: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 2730: 3 -> 10 (AXI_WRITE)\n    inject_packet(3, 10, 64, "AXI_WRITE");\n    // Packet 2731: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 2732: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 2733: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Packet 2734: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 2735: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 573\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 573\n    // Packet 2736: 1 -> 3 (AXI_READ)\n    inject_packet(1, 3, 64, "AXI_READ");\n    // Packet 2737: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 2738: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 2739: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Packet 2740: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 574\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 574\n    // Packet 2741: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 2742: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 2743: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Packet 2744: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Packet 2745: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Packet 2746: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 575\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 575\n    // Packet 2747: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 2748: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 2749: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 2750: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 2751: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 2752: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 2753: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 2754: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 576\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 576\n    // Packet 2755: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 2756: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 2757: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 2758: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 2759: 13 -> 9 (AXI_WRITE)\n    inject_packet(13, 9, 64, "AXI_WRITE");\n    // Wait until cycle 577\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 577\n    // Packet 2760: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 2761: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 2762: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 2763: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Wait until cycle 578\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 578\n    // Packet 2764: 9 -> 7 (AXI_WRITE)\n    inject_packet(9, 7, 64, "AXI_WRITE");\n    // Packet 2765: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Wait until cycle 579\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 579\n    // Packet 2766: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 2767: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 2768: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 2769: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Packet 2770: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 580\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 580\n    // Packet 2771: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 2772: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 2773: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 2774: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 2775: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 2776: 12 -> 3 (AXI_WRITE)\n    inject_packet(12, 3, 64, "AXI_WRITE");\n    // Wait until cycle 581\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 581\n    // Packet 2777: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2778: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 2779: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Packet 2780: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 2781: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 2782: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 2783: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Packet 2784: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 2785: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Packet 2786: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 582\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 582\n    // Packet 2787: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 2788: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 2789: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 2790: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 2791: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 2792: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 2793: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 2794: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 583\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 583\n    // Packet 2795: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 2796: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 2797: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 2798: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Packet 2799: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 584\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 584\n    // Packet 2800: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 2801: 10 -> 4 (AXI_READ)\n    inject_packet(10, 4, 64, "AXI_READ");\n    // Wait until cycle 585\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 585\n    // Packet 2802: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 2803: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 2804: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 2805: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Wait until cycle 586\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 586\n    // Packet 2806: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 2807: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 2808: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 2809: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 2810: 5 -> 15 (AXI_READ)\n    inject_packet(5, 15, 64, "AXI_READ");\n    // Packet 2811: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Packet 2812: 8 -> 1 (AXI_READ)\n    inject_packet(8, 1, 64, "AXI_READ");\n    // Packet 2813: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Wait until cycle 587\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 587\n    // Packet 2814: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 2815: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 2816: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 2817: 8 -> 9 (AXI_READ)\n    inject_packet(8, 9, 64, "AXI_READ");\n    // Packet 2818: 9 -> 0 (AXI_WRITE)\n    inject_packet(9, 0, 64, "AXI_WRITE");\n    // Packet 2819: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Packet 2820: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 588\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 588\n    // Packet 2821: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 2822: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 2823: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 2824: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 2825: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 2826: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Wait until cycle 589\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 589\n    // Packet 2827: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 2828: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Packet 2829: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 590\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 590\n    // Packet 2830: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 2831: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 2832: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Packet 2833: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 2834: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 2835: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 2836: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 591\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 591\n    // Packet 2837: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 2838: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Packet 2839: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 593\n    repeat(2) @(posedge clk);\n    // Inject packets at cycle 593\n    // Packet 2840: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 2841: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 2842: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 2843: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 2844: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 594\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 594\n    // Packet 2845: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 2846: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 2847: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 2848: 5 -> 15 (AXI_READ)\n    inject_packet(5, 15, 64, "AXI_READ");\n    // Packet 2849: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 2850: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Wait until cycle 595\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 595\n    // Packet 2851: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 2852: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 2853: 5 -> 9 (AXI_WRITE)\n    inject_packet(5, 9, 64, "AXI_WRITE");\n    // Packet 2854: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 2855: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Wait until cycle 596\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 596\n    // Packet 2856: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 2857: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Packet 2858: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 597\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 597\n    // Packet 2859: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 2860: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 2861: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 2862: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Wait until cycle 598\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 598\n    // Packet 2863: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 2864: 3 -> 5 (AXI_WRITE)\n    inject_packet(3, 5, 64, "AXI_WRITE");\n    // Packet 2865: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 2866: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 2867: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 599\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 599\n    // Packet 2868: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 2869: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 2870: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 2871: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 2872: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 2873: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Wait until cycle 600\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 600\n    // Packet 2874: 3 -> 8 (AXI_READ)\n    inject_packet(3, 8, 64, "AXI_READ");\n    // Packet 2875: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 2876: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 2877: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 2878: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Packet 2879: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 601\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 601\n    // Packet 2880: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Wait until cycle 602\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 602\n    // Packet 2881: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 2882: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 2883: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Wait until cycle 603\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 603\n    // Packet 2884: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 2885: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Wait until cycle 604\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 604\n    // Packet 2886: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 2887: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Packet 2888: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Wait until cycle 605\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 605\n    // Packet 2889: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 2890: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 2891: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 2892: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 2893: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Wait until cycle 606\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 606\n    // Packet 2894: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 2895: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 2896: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 2897: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 2898: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 2899: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 2900: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Wait until cycle 607\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 607\n    // Packet 2901: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 2902: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 2903: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 2904: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Packet 2905: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 608\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 608\n    // Packet 2906: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 2907: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 2908: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 2909: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 2910: 13 -> 9 (AXI_WRITE)\n    inject_packet(13, 9, 64, "AXI_WRITE");\n    // Wait until cycle 609\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 609\n    // Packet 2911: 0 -> 12 (AXI_READ)\n    inject_packet(0, 12, 64, "AXI_READ");\n    // Packet 2912: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 2913: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Wait until cycle 610\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 610\n    // Packet 2914: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 2915: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 2916: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 2917: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 2918: 12 -> 14 (AXI_READ)\n    inject_packet(12, 14, 64, "AXI_READ");\n    // Packet 2919: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Wait until cycle 611\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 611\n    // Packet 2920: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 2921: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 2922: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 2923: 14 -> 4 (AXI_WRITE)\n    inject_packet(14, 4, 64, "AXI_WRITE");\n    // Wait until cycle 612\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 612\n    // Packet 2924: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 2925: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 2926: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Packet 2927: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 2928: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Packet 2929: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 613\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 613\n    // Packet 2930: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 2931: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 2932: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 2933: 10 -> 3 (AXI_READ)\n    inject_packet(10, 3, 64, "AXI_READ");\n    // Packet 2934: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Packet 2935: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Wait until cycle 614\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 614\n    // Packet 2936: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 2937: 6 -> 2 (AXI_WRITE)\n    inject_packet(6, 2, 64, "AXI_WRITE");\n    // Packet 2938: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 2939: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Packet 2940: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Wait until cycle 615\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 615\n    // Packet 2941: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 2942: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 2943: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 2944: 15 -> 1 (AXI_WRITE)\n    inject_packet(15, 1, 64, "AXI_WRITE");\n    // Wait until cycle 616\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 616\n    // Packet 2945: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 2946: 9 -> 11 (AXI_READ)\n    inject_packet(9, 11, 64, "AXI_READ");\n    // Packet 2947: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Wait until cycle 617\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 617\n    // Packet 2948: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 2949: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 2950: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 2951: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Packet 2952: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 2953: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Packet 2954: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 618\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 618\n    // Packet 2955: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 2956: 7 -> 4 (AXI_WRITE)\n    inject_packet(7, 4, 64, "AXI_WRITE");\n    // Packet 2957: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Packet 2958: 12 -> 9 (AXI_READ)\n    inject_packet(12, 9, 64, "AXI_READ");\n    // Packet 2959: 13 -> 4 (AXI_WRITE)\n    inject_packet(13, 4, 64, "AXI_WRITE");\n    // Wait until cycle 619\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 619\n    // Packet 2960: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 2961: 6 -> 0 (AXI_WRITE)\n    inject_packet(6, 0, 64, "AXI_WRITE");\n    // Packet 2962: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Wait until cycle 620\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 620\n    // Packet 2963: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Wait until cycle 621\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 621\n    // Packet 2964: 1 -> 15 (AXI_READ)\n    inject_packet(1, 15, 64, "AXI_READ");\n    // Packet 2965: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 2966: 3 -> 7 (AXI_READ)\n    inject_packet(3, 7, 64, "AXI_READ");\n    // Packet 2967: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 2968: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 2969: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 2970: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 2971: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 2972: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 2973: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 622\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 622\n    // Packet 2974: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 2975: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 2976: 5 -> 9 (AXI_READ)\n    inject_packet(5, 9, 64, "AXI_READ");\n    // Packet 2977: 7 -> 6 (AXI_WRITE)\n    inject_packet(7, 6, 64, "AXI_WRITE");\n    // Packet 2978: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 2979: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 623\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 623\n    // Packet 2980: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 2981: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 2982: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 2983: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 2984: 5 -> 15 (AXI_READ)\n    inject_packet(5, 15, 64, "AXI_READ");\n    // Packet 2985: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 2986: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 624\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 624\n    // Packet 2987: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 2988: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 2989: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 2990: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 2991: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 2992: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 2993: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 625\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 625\n    // Packet 2994: 2 -> 10 (AXI_READ)\n    inject_packet(2, 10, 64, "AXI_READ");\n    // Packet 2995: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 2996: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 2997: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 626\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 626\n    // Packet 2998: 0 -> 9 (AXI_READ)\n    inject_packet(0, 9, 64, "AXI_READ");\n    // Packet 2999: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 3000: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 3001: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 3002: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 3003: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 3004: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Packet 3005: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Wait until cycle 627\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 627\n    // Packet 3006: 3 -> 2 (AXI_READ)\n    inject_packet(3, 2, 64, "AXI_READ");\n    // Packet 3007: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 3008: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 3009: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 3010: 14 -> 4 (AXI_WRITE)\n    inject_packet(14, 4, 64, "AXI_WRITE");\n    // Packet 3011: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 628\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 628\n    // Packet 3012: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 3013: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 629\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 629\n    // Packet 3014: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 3015: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 3016: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 3017: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 3018: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 630\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 630\n    // Packet 3019: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 3020: 5 -> 0 (AXI_WRITE)\n    inject_packet(5, 0, 64, "AXI_WRITE");\n    // Packet 3021: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 3022: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Wait until cycle 631\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 631\n    // Packet 3023: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 3024: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 3025: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 3026: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 3027: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 632\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 632\n    // Packet 3028: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 3029: 2 -> 5 (AXI_WRITE)\n    inject_packet(2, 5, 64, "AXI_WRITE");\n    // Packet 3030: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 3031: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 3032: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 3033: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 3034: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Wait until cycle 633\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 633\n    // Packet 3035: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 3036: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 3037: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 634\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 634\n    // Packet 3038: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 3039: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 3040: 3 -> 13 (AXI_WRITE)\n    inject_packet(3, 13, 64, "AXI_WRITE");\n    // Packet 3041: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 3042: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 3043: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Wait until cycle 635\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 635\n    // Packet 3044: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 3045: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 3046: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Wait until cycle 636\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 636\n    // Packet 3047: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 3048: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 3049: 10 -> 2 (AXI_READ)\n    inject_packet(10, 2, 64, "AXI_READ");\n    // Packet 3050: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 3051: 14 -> 4 (AXI_READ)\n    inject_packet(14, 4, 64, "AXI_READ");\n    // Wait until cycle 637\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 637\n    // Packet 3052: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 3053: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 3054: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Wait until cycle 638\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 638\n    // Packet 3055: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 3056: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 3057: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 3058: 8 -> 15 (AXI_READ)\n    inject_packet(8, 15, 64, "AXI_READ");\n    // Packet 3059: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 3060: 13 -> 5 (AXI_READ)\n    inject_packet(13, 5, 64, "AXI_READ");\n    // Wait until cycle 639\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 639\n    // Packet 3061: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 3062: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 3063: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 3064: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Wait until cycle 640\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 640\n    // Packet 3065: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 3066: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 3067: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 3068: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 3069: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 3070: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 3071: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 641\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 641\n    // Packet 3072: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 3073: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 3074: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 3075: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 3076: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 642\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 642\n    // Packet 3077: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Wait until cycle 643\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 643\n    // Packet 3078: 1 -> 9 (AXI_WRITE)\n    inject_packet(1, 9, 64, "AXI_WRITE");\n    // Packet 3079: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 3080: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 3081: 7 -> 13 (AXI_WRITE)\n    inject_packet(7, 13, 64, "AXI_WRITE");\n    // Packet 3082: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Packet 3083: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 644\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 644\n    // Packet 3084: 7 -> 13 (AXI_WRITE)\n    inject_packet(7, 13, 64, "AXI_WRITE");\n    // Packet 3085: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 3086: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 645\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 645\n    // Packet 3087: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 3088: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 3089: 14 -> 9 (AXI_WRITE)\n    inject_packet(14, 9, 64, "AXI_WRITE");\n    // Wait until cycle 646\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 646\n    // Packet 3090: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 3091: 1 -> 9 (AXI_WRITE)\n    inject_packet(1, 9, 64, "AXI_WRITE");\n    // Packet 3092: 6 -> 9 (AXI_WRITE)\n    inject_packet(6, 9, 64, "AXI_WRITE");\n    // Packet 3093: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Packet 3094: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Wait until cycle 647\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 647\n    // Packet 3095: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 3096: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 3097: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 3098: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 3099: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Packet 3100: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Wait until cycle 648\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 648\n    // Packet 3101: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 3102: 6 -> 4 (AXI_READ)\n    inject_packet(6, 4, 64, "AXI_READ");\n    // Wait until cycle 649\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 649\n    // Packet 3103: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 3104: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 3105: 7 -> 8 (AXI_READ)\n    inject_packet(7, 8, 64, "AXI_READ");\n    // Packet 3106: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 3107: 12 -> 13 (AXI_READ)\n    inject_packet(12, 13, 64, "AXI_READ");\n    // Wait until cycle 650\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 650\n    // Packet 3108: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 3109: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 3110: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 3111: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 3112: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 3113: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Packet 3114: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 651\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 651\n    // Packet 3115: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 3116: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 3117: 10 -> 7 (AXI_READ)\n    inject_packet(10, 7, 64, "AXI_READ");\n    // Wait until cycle 652\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 652\n    // Packet 3118: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 3119: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 3120: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 3121: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Wait until cycle 653\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 653\n    // Packet 3122: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 3123: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 3124: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 3125: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 654\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 654\n    // Packet 3126: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 3127: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 655\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 655\n    // Packet 3128: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 3129: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 3130: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 3131: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 3132: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 3133: 10 -> 5 (AXI_WRITE)\n    inject_packet(10, 5, 64, "AXI_WRITE");\n    // Packet 3134: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Packet 3135: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 656\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 656\n    // Packet 3136: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 3137: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 3138: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 3139: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Wait until cycle 657\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 657\n    // Packet 3140: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 3141: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 3142: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Packet 3143: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Packet 3144: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 658\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 658\n    // Packet 3145: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Packet 3146: 5 -> 13 (AXI_READ)\n    inject_packet(5, 13, 64, "AXI_READ");\n    // Packet 3147: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 3148: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 3149: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Wait until cycle 659\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 659\n    // Packet 3150: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Wait until cycle 660\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 660\n    // Packet 3151: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 3152: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 3153: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 3154: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 3155: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Wait until cycle 661\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 661\n    // Packet 3156: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 3157: 4 -> 1 (AXI_WRITE)\n    inject_packet(4, 1, 64, "AXI_WRITE");\n    // Packet 3158: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 3159: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 3160: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 3161: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Packet 3162: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Wait until cycle 662\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 662\n    // Packet 3163: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 3164: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 3165: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 3166: 8 -> 4 (AXI_READ)\n    inject_packet(8, 4, 64, "AXI_READ");\n    // Packet 3167: 12 -> 14 (AXI_READ)\n    inject_packet(12, 14, 64, "AXI_READ");\n    // Packet 3168: 15 -> 3 (AXI_WRITE)\n    inject_packet(15, 3, 64, "AXI_WRITE");\n    // Wait until cycle 663\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 663\n    // Packet 3169: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 3170: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 3171: 8 -> 12 (AXI_READ)\n    inject_packet(8, 12, 64, "AXI_READ");\n    // Packet 3172: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 664\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 664\n    // Packet 3173: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 3174: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 3175: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 3176: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 3177: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 3178: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Packet 3179: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 665\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 665\n    // Packet 3180: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Packet 3181: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 666\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 666\n    // Packet 3182: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 3183: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 3184: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Packet 3185: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 667\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 667\n    // Packet 3186: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 3187: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 3188: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 3189: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 3190: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 3191: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 3192: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Wait until cycle 668\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 668\n    // Packet 3193: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 3194: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 3195: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Packet 3196: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Packet 3197: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 669\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 669\n    // Packet 3198: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 3199: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 3200: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 3201: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Wait until cycle 670\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 670\n    // Packet 3202: 1 -> 3 (AXI_WRITE)\n    inject_packet(1, 3, 64, "AXI_WRITE");\n    // Wait until cycle 671\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 671\n    // Packet 3203: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 3204: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 3205: 9 -> 13 (AXI_READ)\n    inject_packet(9, 13, 64, "AXI_READ");\n    // Wait until cycle 672\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 672\n    // Packet 3206: 0 -> 10 (AXI_READ)\n    inject_packet(0, 10, 64, "AXI_READ");\n    // Packet 3207: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 3208: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 3209: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 673\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 673\n    // Packet 3210: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 3211: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Packet 3212: 6 -> 0 (AXI_WRITE)\n    inject_packet(6, 0, 64, "AXI_WRITE");\n    // Packet 3213: 7 -> 4 (AXI_WRITE)\n    inject_packet(7, 4, 64, "AXI_WRITE");\n    // Packet 3214: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 3215: 11 -> 9 (AXI_READ)\n    inject_packet(11, 9, 64, "AXI_READ");\n    // Packet 3216: 13 -> 5 (AXI_READ)\n    inject_packet(13, 5, 64, "AXI_READ");\n    // Wait until cycle 674\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 674\n    // Packet 3217: 3 -> 12 (AXI_WRITE)\n    inject_packet(3, 12, 64, "AXI_WRITE");\n    // Packet 3218: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 3219: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 3220: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 3221: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 3222: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Wait until cycle 675\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 675\n    // Packet 3223: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 3224: 15 -> 0 (AXI_WRITE)\n    inject_packet(15, 0, 64, "AXI_WRITE");\n    // Wait until cycle 676\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 676\n    // Packet 3225: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 3226: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 3227: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 3228: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 3229: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Wait until cycle 677\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 677\n    // Packet 3230: 1 -> 10 (AXI_READ)\n    inject_packet(1, 10, 64, "AXI_READ");\n    // Packet 3231: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 3232: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 3233: 10 -> 2 (AXI_READ)\n    inject_packet(10, 2, 64, "AXI_READ");\n    // Wait until cycle 678\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 678\n    // Packet 3234: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 3235: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 3236: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 3237: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 3238: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 3239: 11 -> 9 (AXI_READ)\n    inject_packet(11, 9, 64, "AXI_READ");\n    // Wait until cycle 679\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 679\n    // Packet 3240: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 3241: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 3242: 6 -> 9 (AXI_WRITE)\n    inject_packet(6, 9, 64, "AXI_WRITE");\n    // Packet 3243: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 3244: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 3245: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Wait until cycle 680\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 680\n    // Packet 3246: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 3247: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 3248: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 3249: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 3250: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Wait until cycle 681\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 681\n    // Packet 3251: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 3252: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 3253: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 3254: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 3255: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 3256: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 3257: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 3258: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Wait until cycle 682\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 682\n    // Packet 3259: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 3260: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 3261: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 3262: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 3263: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 683\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 683\n    // Packet 3264: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 3265: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 3266: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 3267: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 3268: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 3269: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Wait until cycle 684\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 684\n    // Packet 3270: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 3271: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 3272: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 3273: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Packet 3274: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 685\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 685\n    // Packet 3275: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 3276: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 3277: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 3278: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 686\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 686\n    // Packet 3279: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 3280: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 3281: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 3282: 14 -> 9 (AXI_WRITE)\n    inject_packet(14, 9, 64, "AXI_WRITE");\n    // Wait until cycle 687\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 687\n    // Packet 3283: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 3284: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 3285: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 3286: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Packet 3287: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Wait until cycle 688\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 688\n    // Packet 3288: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 3289: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 3290: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Packet 3291: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 689\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 689\n    // Packet 3292: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 3293: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Packet 3294: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 3295: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 3296: 13 -> 1 (AXI_WRITE)\n    inject_packet(13, 1, 64, "AXI_WRITE");\n    // Packet 3297: 14 -> 2 (AXI_READ)\n    inject_packet(14, 2, 64, "AXI_READ");\n    // Wait until cycle 690\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 690\n    // Packet 3298: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 3299: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 3300: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Wait until cycle 691\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 691\n    // Packet 3301: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 3302: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 3303: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 692\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 692\n    // Packet 3304: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 3305: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 3306: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 3307: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Wait until cycle 693\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 693\n    // Packet 3308: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 3309: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 3310: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 3311: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 3312: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Packet 3313: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 694\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 694\n    // Packet 3314: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 3315: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 3316: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 3317: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 3318: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Packet 3319: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Wait until cycle 695\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 695\n    // Packet 3320: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 3321: 2 -> 11 (AXI_WRITE)\n    inject_packet(2, 11, 64, "AXI_WRITE");\n    // Packet 3322: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 3323: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 3324: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 3325: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Wait until cycle 696\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 696\n    // Packet 3326: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 3327: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 3328: 12 -> 3 (AXI_WRITE)\n    inject_packet(12, 3, 64, "AXI_WRITE");\n    // Wait until cycle 697\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 697\n    // Packet 3329: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 3330: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 3331: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 3332: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 698\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 698\n    // Packet 3333: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 3334: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 3335: 8 -> 9 (AXI_READ)\n    inject_packet(8, 9, 64, "AXI_READ");\n    // Packet 3336: 12 -> 1 (AXI_WRITE)\n    inject_packet(12, 1, 64, "AXI_WRITE");\n    // Packet 3337: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Wait until cycle 699\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 699\n    // Packet 3338: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Wait until cycle 700\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 700\n    // Packet 3339: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 3340: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 3341: 9 -> 15 (AXI_WRITE)\n    inject_packet(9, 15, 64, "AXI_WRITE");\n    // Packet 3342: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 3343: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 701\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 701\n    // Packet 3344: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 3345: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 3346: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 3347: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 3348: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 3349: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Wait until cycle 702\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 702\n    // Packet 3350: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 3351: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 3352: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Packet 3353: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Packet 3354: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Wait until cycle 703\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 703\n    // Packet 3355: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 3356: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 3357: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 3358: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 3359: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Wait until cycle 704\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 704\n    // Packet 3360: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 3361: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 3362: 10 -> 13 (AXI_READ)\n    inject_packet(10, 13, 64, "AXI_READ");\n    // Packet 3363: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 3364: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 705\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 705\n    // Packet 3365: 6 -> 2 (AXI_WRITE)\n    inject_packet(6, 2, 64, "AXI_WRITE");\n    // Packet 3366: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 3367: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 3368: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Wait until cycle 706\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 706\n    // Packet 3369: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 3370: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 3371: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 707\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 707\n    // Packet 3372: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 3373: 1 -> 8 (AXI_WRITE)\n    inject_packet(1, 8, 64, "AXI_WRITE");\n    // Packet 3374: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 3375: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 3376: 7 -> 9 (AXI_WRITE)\n    inject_packet(7, 9, 64, "AXI_WRITE");\n    // Packet 3377: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Packet 3378: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 3379: 15 -> 13 (AXI_WRITE)\n    inject_packet(15, 13, 64, "AXI_WRITE");\n    // Wait until cycle 708\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 708\n    // Packet 3380: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 3381: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 3382: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 3383: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 3384: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 709\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 709\n    // Packet 3385: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 3386: 1 -> 15 (AXI_READ)\n    inject_packet(1, 15, 64, "AXI_READ");\n    // Packet 3387: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Packet 3388: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 3389: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 3390: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Wait until cycle 710\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 710\n    // Packet 3391: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 3392: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 3393: 6 -> 8 (AXI_WRITE)\n    inject_packet(6, 8, 64, "AXI_WRITE");\n    // Packet 3394: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 711\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 711\n    // Packet 3395: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 3396: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 3397: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 712\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 712\n    // Packet 3398: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 3399: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 3400: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 3401: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 3402: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 3403: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Packet 3404: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 713\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 713\n    // Packet 3405: 2 -> 0 (AXI_WRITE)\n    inject_packet(2, 0, 64, "AXI_WRITE");\n    // Packet 3406: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 3407: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 3408: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 3409: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 3410: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Packet 3411: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Packet 3412: 14 -> 4 (AXI_WRITE)\n    inject_packet(14, 4, 64, "AXI_WRITE");\n    // Wait until cycle 714\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 714\n    // Packet 3413: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 3414: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 3415: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 715\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 715\n    // Packet 3416: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 3417: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 3418: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 3419: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 3420: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Wait until cycle 716\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 716\n    // Packet 3421: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 3422: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 3423: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 3424: 13 -> 0 (AXI_WRITE)\n    inject_packet(13, 0, 64, "AXI_WRITE");\n    // Wait until cycle 717\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 717\n    // Packet 3425: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 3426: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Wait until cycle 718\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 718\n    // Packet 3427: 0 -> 14 (AXI_READ)\n    inject_packet(0, 14, 64, "AXI_READ");\n    // Packet 3428: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 3429: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 3430: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 719\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 719\n    // Packet 3431: 2 -> 1 (AXI_WRITE)\n    inject_packet(2, 1, 64, "AXI_WRITE");\n    // Packet 3432: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 3433: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Packet 3434: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 720\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 720\n    // Packet 3435: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 3436: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 3437: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 3438: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 3439: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 3440: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 3441: 13 -> 2 (AXI_WRITE)\n    inject_packet(13, 2, 64, "AXI_WRITE");\n    // Wait until cycle 721\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 721\n    // Packet 3442: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 3443: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 3444: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 3445: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 3446: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 3447: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Wait until cycle 722\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 722\n    // Packet 3448: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 3449: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 3450: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 3451: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 723\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 723\n    // Packet 3452: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 3453: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Wait until cycle 724\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 724\n    // Packet 3454: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 3455: 4 -> 8 (AXI_READ)\n    inject_packet(4, 8, 64, "AXI_READ");\n    // Packet 3456: 10 -> 7 (AXI_READ)\n    inject_packet(10, 7, 64, "AXI_READ");\n    // Packet 3457: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Packet 3458: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Packet 3459: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 725\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 725\n    // Packet 3460: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 3461: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 3462: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 3463: 8 -> 14 (AXI_WRITE)\n    inject_packet(8, 14, 64, "AXI_WRITE");\n    // Packet 3464: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 726\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 726\n    // Packet 3465: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 3466: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 3467: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Wait until cycle 727\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 727\n    // Packet 3468: 1 -> 3 (AXI_READ)\n    inject_packet(1, 3, 64, "AXI_READ");\n    // Packet 3469: 6 -> 8 (AXI_WRITE)\n    inject_packet(6, 8, 64, "AXI_WRITE");\n    // Packet 3470: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Wait until cycle 728\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 728\n    // Packet 3471: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 3472: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 3473: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Wait until cycle 729\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 729\n    // Packet 3474: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 3475: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 3476: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Wait until cycle 730\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 730\n    // Packet 3477: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 3478: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 3479: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Packet 3480: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 731\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 731\n    // Packet 3481: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 3482: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 3483: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Wait until cycle 732\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 732\n    // Packet 3484: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 3485: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 3486: 9 -> 0 (AXI_WRITE)\n    inject_packet(9, 0, 64, "AXI_WRITE");\n    // Wait until cycle 733\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 733\n    // Packet 3487: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 3488: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 3489: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 3490: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Packet 3491: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Wait until cycle 734\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 734\n    // Packet 3492: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 3493: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 3494: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 3495: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 3496: 9 -> 0 (AXI_READ)\n    inject_packet(9, 0, 64, "AXI_READ");\n    // Packet 3497: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Packet 3498: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 735\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 735\n    // Packet 3499: 4 -> 3 (AXI_READ)\n    inject_packet(4, 3, 64, "AXI_READ");\n    // Packet 3500: 9 -> 0 (AXI_READ)\n    inject_packet(9, 0, 64, "AXI_READ");\n    // Packet 3501: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 3502: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 736\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 736\n    // Packet 3503: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Packet 3504: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Wait until cycle 737\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 737\n    // Packet 3505: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 3506: 3 -> 5 (AXI_WRITE)\n    inject_packet(3, 5, 64, "AXI_WRITE");\n    // Packet 3507: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 3508: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Packet 3509: 10 -> 13 (AXI_READ)\n    inject_packet(10, 13, 64, "AXI_READ");\n    // Packet 3510: 11 -> 6 (AXI_READ)\n    inject_packet(11, 6, 64, "AXI_READ");\n    // Packet 3511: 12 -> 13 (AXI_READ)\n    inject_packet(12, 13, 64, "AXI_READ");\n    // Packet 3512: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 738\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 738\n    // Packet 3513: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 3514: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 3515: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Wait until cycle 739\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 739\n    // Packet 3516: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 3517: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Wait until cycle 740\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 740\n    // Packet 3518: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 3519: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 3520: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 3521: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 3522: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 3523: 14 -> 5 (AXI_READ)\n    inject_packet(14, 5, 64, "AXI_READ");\n    // Wait until cycle 741\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 741\n    // Packet 3524: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 3525: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 3526: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 3527: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 3528: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 3529: 12 -> 13 (AXI_READ)\n    inject_packet(12, 13, 64, "AXI_READ");\n    // Wait until cycle 742\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 742\n    // Packet 3530: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 3531: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 3532: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 3533: 10 -> 1 (AXI_READ)\n    inject_packet(10, 1, 64, "AXI_READ");\n    // Packet 3534: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Wait until cycle 743\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 743\n    // Packet 3535: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 3536: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 3537: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 3538: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Packet 3539: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 3540: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Wait until cycle 744\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 744\n    // Packet 3541: 7 -> 9 (AXI_WRITE)\n    inject_packet(7, 9, 64, "AXI_WRITE");\n    // Packet 3542: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 3543: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Wait until cycle 745\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 745\n    // Packet 3544: 1 -> 4 (AXI_WRITE)\n    inject_packet(1, 4, 64, "AXI_WRITE");\n    // Packet 3545: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 3546: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 3547: 11 -> 6 (AXI_READ)\n    inject_packet(11, 6, 64, "AXI_READ");\n    // Wait until cycle 746\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 746\n    // Packet 3548: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 3549: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Wait until cycle 747\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 747\n    // Packet 3550: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 3551: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 3552: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 3553: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 3554: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Wait until cycle 748\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 748\n    // Packet 3555: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Wait until cycle 749\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 749\n    // Packet 3556: 1 -> 4 (AXI_WRITE)\n    inject_packet(1, 4, 64, "AXI_WRITE");\n    // Packet 3557: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 3558: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Packet 3559: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 750\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 750\n    // Packet 3560: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 3561: 10 -> 14 (AXI_READ)\n    inject_packet(10, 14, 64, "AXI_READ");\n    // Packet 3562: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 3563: 12 -> 5 (AXI_READ)\n    inject_packet(12, 5, 64, "AXI_READ");\n    // Packet 3564: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 3565: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 751\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 751\n    // Packet 3566: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 3567: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 3568: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 3569: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 3570: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Wait until cycle 752\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 752\n    // Packet 3571: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 3572: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 3573: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 3574: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 3575: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 3576: 7 -> 14 (AXI_WRITE)\n    inject_packet(7, 14, 64, "AXI_WRITE");\n    // Packet 3577: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 3578: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 3579: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 753\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 753\n    // Packet 3580: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 3581: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 3582: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 3583: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 3584: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 3585: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 754\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 754\n    // Packet 3586: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 3587: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 3588: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 3589: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 3590: 11 -> 0 (AXI_READ)\n    inject_packet(11, 0, 64, "AXI_READ");\n    // Packet 3591: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Packet 3592: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Packet 3593: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 755\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 755\n    // Packet 3594: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 3595: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 3596: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Packet 3597: 11 -> 9 (AXI_READ)\n    inject_packet(11, 9, 64, "AXI_READ");\n    // Packet 3598: 14 -> 4 (AXI_WRITE)\n    inject_packet(14, 4, 64, "AXI_WRITE");\n    // Wait until cycle 756\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 756\n    // Packet 3599: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 3600: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 3601: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 3602: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 3603: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 3604: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Packet 3605: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 3606: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 758\n    repeat(2) @(posedge clk);\n    // Inject packets at cycle 758\n    // Packet 3607: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 3608: 1 -> 8 (AXI_WRITE)\n    inject_packet(1, 8, 64, "AXI_WRITE");\n    // Packet 3609: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 3610: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 3611: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 3612: 12 -> 14 (AXI_READ)\n    inject_packet(12, 14, 64, "AXI_READ");\n    // Packet 3613: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Packet 3614: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Packet 3615: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 759\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 759\n    // Packet 3616: 1 -> 15 (AXI_WRITE)\n    inject_packet(1, 15, 64, "AXI_WRITE");\n    // Packet 3617: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 3618: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 3619: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 3620: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 3621: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 3622: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Packet 3623: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 3624: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 760\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 760\n    // Packet 3625: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 3626: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 3627: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 3628: 13 -> 9 (AXI_WRITE)\n    inject_packet(13, 9, 64, "AXI_WRITE");\n    // Packet 3629: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 761\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 761\n    // Packet 3630: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 3631: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 3632: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Packet 3633: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Packet 3634: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 762\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 762\n    // Packet 3635: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 3636: 12 -> 9 (AXI_READ)\n    inject_packet(12, 9, 64, "AXI_READ");\n    // Packet 3637: 13 -> 10 (AXI_WRITE)\n    inject_packet(13, 10, 64, "AXI_WRITE");\n    // Packet 3638: 15 -> 5 (AXI_WRITE)\n    inject_packet(15, 5, 64, "AXI_WRITE");\n    // Wait until cycle 763\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 763\n    // Packet 3639: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 3640: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 3641: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Packet 3642: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 3643: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Packet 3644: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Wait until cycle 764\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 764\n    // Packet 3645: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 3646: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 3647: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 3648: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Wait until cycle 765\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 765\n    // Packet 3649: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 3650: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 3651: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 3652: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Packet 3653: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Packet 3654: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 766\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 766\n    // Packet 3655: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 3656: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 3657: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Wait until cycle 767\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 767\n    // Packet 3658: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 3659: 5 -> 3 (AXI_WRITE)\n    inject_packet(5, 3, 64, "AXI_WRITE");\n    // Packet 3660: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 3661: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Packet 3662: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Packet 3663: 14 -> 15 (AXI_WRITE)\n    inject_packet(14, 15, 64, "AXI_WRITE");\n    // Wait until cycle 768\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 768\n    // Packet 3664: 0 -> 9 (AXI_READ)\n    inject_packet(0, 9, 64, "AXI_READ");\n    // Packet 3665: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 3666: 3 -> 12 (AXI_WRITE)\n    inject_packet(3, 12, 64, "AXI_WRITE");\n    // Packet 3667: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 3668: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 3669: 11 -> 2 (AXI_READ)\n    inject_packet(11, 2, 64, "AXI_READ");\n    // Wait until cycle 769\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 769\n    // Packet 3670: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 3671: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 3672: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 3673: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Packet 3674: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Packet 3675: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 770\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 770\n    // Packet 3676: 0 -> 14 (AXI_WRITE)\n    inject_packet(0, 14, 64, "AXI_WRITE");\n    // Packet 3677: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 3678: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Packet 3679: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 771\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 771\n    // Packet 3680: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 3681: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 3682: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 3683: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 3684: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 3685: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Wait until cycle 772\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 772\n    // Packet 3686: 6 -> 9 (AXI_WRITE)\n    inject_packet(6, 9, 64, "AXI_WRITE");\n    // Packet 3687: 10 -> 13 (AXI_READ)\n    inject_packet(10, 13, 64, "AXI_READ");\n    // Packet 3688: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Packet 3689: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 773\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 773\n    // Packet 3690: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 3691: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 3692: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 3693: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 3694: 11 -> 3 (AXI_READ)\n    inject_packet(11, 3, 64, "AXI_READ");\n    // Packet 3695: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Packet 3696: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 774\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 774\n    // Packet 3697: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 3698: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 3699: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 3700: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 3701: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 3702: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 3703: 14 -> 4 (AXI_WRITE)\n    inject_packet(14, 4, 64, "AXI_WRITE");\n    // Packet 3704: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 775\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 775\n    // Packet 3705: 3 -> 8 (AXI_READ)\n    inject_packet(3, 8, 64, "AXI_READ");\n    // Packet 3706: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 3707: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 3708: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Wait until cycle 776\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 776\n    // Packet 3709: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 3710: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 3711: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Wait until cycle 777\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 777\n    // Packet 3712: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 3713: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 3714: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 3715: 8 -> 2 (AXI_WRITE)\n    inject_packet(8, 2, 64, "AXI_WRITE");\n    // Packet 3716: 15 -> 4 (AXI_READ)\n    inject_packet(15, 4, 64, "AXI_READ");\n    // Wait until cycle 778\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 778\n    // Packet 3717: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 3718: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 3719: 7 -> 8 (AXI_READ)\n    inject_packet(7, 8, 64, "AXI_READ");\n    // Packet 3720: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 3721: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 3722: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Packet 3723: 14 -> 0 (AXI_READ)\n    inject_packet(14, 0, 64, "AXI_READ");\n    // Wait until cycle 779\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 779\n    // Packet 3724: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 3725: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 3726: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 3727: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 3728: 12 -> 0 (AXI_WRITE)\n    inject_packet(12, 0, 64, "AXI_WRITE");\n    // Packet 3729: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Packet 3730: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 780\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 780\n    // Packet 3731: 1 -> 15 (AXI_WRITE)\n    inject_packet(1, 15, 64, "AXI_WRITE");\n    // Packet 3732: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 3733: 6 -> 4 (AXI_WRITE)\n    inject_packet(6, 4, 64, "AXI_WRITE");\n    // Packet 3734: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 781\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 781\n    // Packet 3735: 1 -> 6 (AXI_WRITE)\n    inject_packet(1, 6, 64, "AXI_WRITE");\n    // Packet 3736: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 3737: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 3738: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Packet 3739: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Wait until cycle 782\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 782\n    // Packet 3740: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 3741: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 3742: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 3743: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 3744: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 3745: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 3746: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Packet 3747: 11 -> 3 (AXI_WRITE)\n    inject_packet(11, 3, 64, "AXI_WRITE");\n    // Packet 3748: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 783\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 783\n    // Packet 3749: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 3750: 4 -> 9 (AXI_READ)\n    inject_packet(4, 9, 64, "AXI_READ");\n    // Packet 3751: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 3752: 8 -> 9 (AXI_READ)\n    inject_packet(8, 9, 64, "AXI_READ");\n    // Packet 3753: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 3754: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Packet 3755: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 3756: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Wait until cycle 784\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 784\n    // Packet 3757: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 3758: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 3759: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 3760: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 3761: 15 -> 6 (AXI_READ)\n    inject_packet(15, 6, 64, "AXI_READ");\n    // Wait until cycle 785\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 785\n    // Packet 3762: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 3763: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 3764: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 3765: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 3766: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 786\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 786\n    // Packet 3767: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 3768: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 3769: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 3770: 5 -> 12 (AXI_WRITE)\n    inject_packet(5, 12, 64, "AXI_WRITE");\n    // Packet 3771: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 3772: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Wait until cycle 787\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 787\n    // Packet 3773: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Packet 3774: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 3775: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 3776: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 3777: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 3778: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Wait until cycle 788\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 788\n    // Packet 3779: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 3780: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 3781: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 3782: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 3783: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Wait until cycle 789\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 789\n    // Packet 3784: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 3785: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Packet 3786: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Wait until cycle 790\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 790\n    // Packet 3787: 0 -> 2 (AXI_READ)\n    inject_packet(0, 2, 64, "AXI_READ");\n    // Packet 3788: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 3789: 2 -> 4 (AXI_READ)\n    inject_packet(2, 4, 64, "AXI_READ");\n    // Packet 3790: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 3791: 5 -> 12 (AXI_READ)\n    inject_packet(5, 12, 64, "AXI_READ");\n    // Packet 3792: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 791\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 791\n    // Packet 3793: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 3794: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 3795: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 3796: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 792\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 792\n    // Packet 3797: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 3798: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Wait until cycle 793\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 793\n    // Packet 3799: 2 -> 5 (AXI_WRITE)\n    inject_packet(2, 5, 64, "AXI_WRITE");\n    // Packet 3800: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 3801: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Wait until cycle 794\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 794\n    // Packet 3802: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 3803: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 3804: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 3805: 10 -> 7 (AXI_READ)\n    inject_packet(10, 7, 64, "AXI_READ");\n    // Packet 3806: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Packet 3807: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 3808: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Packet 3809: 15 -> 5 (AXI_READ)\n    inject_packet(15, 5, 64, "AXI_READ");\n    // Wait until cycle 795\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 795\n    // Packet 3810: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 3811: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 3812: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 3813: 6 -> 7 (AXI_WRITE)\n    inject_packet(6, 7, 64, "AXI_WRITE");\n    // Packet 3814: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 3815: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 3816: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Wait until cycle 796\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 796\n    // Packet 3817: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Packet 3818: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 3819: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 797\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 797\n    // Packet 3820: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 3821: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 3822: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Wait until cycle 798\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 798\n    // Packet 3823: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 3824: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 3825: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 3826: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 3827: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 3828: 12 -> 5 (AXI_WRITE)\n    inject_packet(12, 5, 64, "AXI_WRITE");\n    // Wait until cycle 799\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 799\n    // Packet 3829: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 3830: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 3831: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 3832: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 3833: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Packet 3834: 13 -> 7 (AXI_WRITE)\n    inject_packet(13, 7, 64, "AXI_WRITE");\n    // Wait until cycle 800\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 800\n    // Packet 3835: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 3836: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 3837: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Packet 3838: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Packet 3839: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 801\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 801\n    // Packet 3840: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 3841: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 3842: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 3843: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 3844: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Packet 3845: 13 -> 14 (AXI_WRITE)\n    inject_packet(13, 14, 64, "AXI_WRITE");\n    // Packet 3846: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Packet 3847: 15 -> 1 (AXI_WRITE)\n    inject_packet(15, 1, 64, "AXI_WRITE");\n    // Wait until cycle 802\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 802\n    // Packet 3848: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 3849: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 3850: 9 -> 3 (AXI_WRITE)\n    inject_packet(9, 3, 64, "AXI_WRITE");\n    // Packet 3851: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 3852: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Packet 3853: 14 -> 9 (AXI_WRITE)\n    inject_packet(14, 9, 64, "AXI_WRITE");\n    // Wait until cycle 803\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 803\n    // Packet 3854: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 3855: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 3856: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 3857: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 3858: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 804\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 804\n    // Packet 3859: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 3860: 5 -> 4 (AXI_WRITE)\n    inject_packet(5, 4, 64, "AXI_WRITE");\n    // Packet 3861: 6 -> 11 (AXI_READ)\n    inject_packet(6, 11, 64, "AXI_READ");\n    // Packet 3862: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 3863: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 3864: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 805\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 805\n    // Packet 3865: 2 -> 5 (AXI_WRITE)\n    inject_packet(2, 5, 64, "AXI_WRITE");\n    // Packet 3866: 7 -> 13 (AXI_WRITE)\n    inject_packet(7, 13, 64, "AXI_WRITE");\n    // Packet 3867: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 3868: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Wait until cycle 806\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 806\n    // Packet 3869: 6 -> 9 (AXI_WRITE)\n    inject_packet(6, 9, 64, "AXI_WRITE");\n    // Packet 3870: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 3871: 11 -> 12 (AXI_READ)\n    inject_packet(11, 12, 64, "AXI_READ");\n    // Wait until cycle 807\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 807\n    // Packet 3872: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 3873: 1 -> 9 (AXI_WRITE)\n    inject_packet(1, 9, 64, "AXI_WRITE");\n    // Packet 3874: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Wait until cycle 808\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 808\n    // Packet 3875: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 3876: 11 -> 8 (AXI_READ)\n    inject_packet(11, 8, 64, "AXI_READ");\n    // Packet 3877: 15 -> 0 (AXI_WRITE)\n    inject_packet(15, 0, 64, "AXI_WRITE");\n    // Wait until cycle 809\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 809\n    // Packet 3878: 3 -> 6 (AXI_READ)\n    inject_packet(3, 6, 64, "AXI_READ");\n    // Packet 3879: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 3880: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Packet 3881: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 3882: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 810\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 810\n    // Packet 3883: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 3884: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 3885: 11 -> 14 (AXI_WRITE)\n    inject_packet(11, 14, 64, "AXI_WRITE");\n    // Packet 3886: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Packet 3887: 15 -> 13 (AXI_WRITE)\n    inject_packet(15, 13, 64, "AXI_WRITE");\n    // Wait until cycle 811\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 811\n    // Packet 3888: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 3889: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 3890: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 3891: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Packet 3892: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 3893: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Packet 3894: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Packet 3895: 15 -> 0 (AXI_WRITE)\n    inject_packet(15, 0, 64, "AXI_WRITE");\n    // Wait until cycle 812\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 812\n    // Packet 3896: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 3897: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 3898: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 3899: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 3900: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 3901: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Packet 3902: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 813\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 813\n    // Packet 3903: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Packet 3904: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 814\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 814\n    // Packet 3905: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 3906: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 3907: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 3908: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 3909: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Packet 3910: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Packet 3911: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 815\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 815\n    // Packet 3912: 8 -> 14 (AXI_WRITE)\n    inject_packet(8, 14, 64, "AXI_WRITE");\n    // Packet 3913: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 3914: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 3915: 11 -> 3 (AXI_READ)\n    inject_packet(11, 3, 64, "AXI_READ");\n    // Packet 3916: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 3917: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 3918: 14 -> 4 (AXI_WRITE)\n    inject_packet(14, 4, 64, "AXI_WRITE");\n    // Wait until cycle 816\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 816\n    // Packet 3919: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 3920: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 3921: 10 -> 8 (AXI_WRITE)\n    inject_packet(10, 8, 64, "AXI_WRITE");\n    // Wait until cycle 817\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 817\n    // Packet 3922: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 3923: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 3924: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 3925: 15 -> 4 (AXI_READ)\n    inject_packet(15, 4, 64, "AXI_READ");\n    // Wait until cycle 818\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 818\n    // Packet 3926: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 3927: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 3928: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 3929: 15 -> 5 (AXI_READ)\n    inject_packet(15, 5, 64, "AXI_READ");\n    // Wait until cycle 819\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 819\n    // Packet 3930: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 3931: 9 -> 14 (AXI_READ)\n    inject_packet(9, 14, 64, "AXI_READ");\n    // Packet 3932: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 3933: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 820\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 820\n    // Packet 3934: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 3935: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 3936: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 3937: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 3938: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 3939: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 3940: 10 -> 12 (AXI_WRITE)\n    inject_packet(10, 12, 64, "AXI_WRITE");\n    // Packet 3941: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 3942: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Packet 3943: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 821\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 821\n    // Packet 3944: 1 -> 0 (AXI_WRITE)\n    inject_packet(1, 0, 64, "AXI_WRITE");\n    // Packet 3945: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 3946: 8 -> 4 (AXI_WRITE)\n    inject_packet(8, 4, 64, "AXI_WRITE");\n    // Packet 3947: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 3948: 11 -> 0 (AXI_READ)\n    inject_packet(11, 0, 64, "AXI_READ");\n    // Packet 3949: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 822\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 822\n    // Packet 3950: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 3951: 5 -> 6 (AXI_READ)\n    inject_packet(5, 6, 64, "AXI_READ");\n    // Packet 3952: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 3953: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 3954: 12 -> 13 (AXI_READ)\n    inject_packet(12, 13, 64, "AXI_READ");\n    // Packet 3955: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Packet 3956: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 823\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 823\n    // Packet 3957: 1 -> 2 (AXI_READ)\n    inject_packet(1, 2, 64, "AXI_READ");\n    // Packet 3958: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 3959: 6 -> 7 (AXI_WRITE)\n    inject_packet(6, 7, 64, "AXI_WRITE");\n    // Packet 3960: 7 -> 1 (AXI_READ)\n    inject_packet(7, 1, 64, "AXI_READ");\n    // Packet 3961: 9 -> 14 (AXI_WRITE)\n    inject_packet(9, 14, 64, "AXI_WRITE");\n    // Packet 3962: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 3963: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 824\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 824\n    // Packet 3964: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 3965: 3 -> 13 (AXI_READ)\n    inject_packet(3, 13, 64, "AXI_READ");\n    // Packet 3966: 4 -> 2 (AXI_READ)\n    inject_packet(4, 2, 64, "AXI_READ");\n    // Packet 3967: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 3968: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 3969: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 3970: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 825\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 825\n    // Packet 3971: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 3972: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 3973: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 3974: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 3975: 8 -> 5 (AXI_WRITE)\n    inject_packet(8, 5, 64, "AXI_WRITE");\n    // Packet 3976: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Wait until cycle 826\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 826\n    // Packet 3977: 1 -> 7 (AXI_WRITE)\n    inject_packet(1, 7, 64, "AXI_WRITE");\n    // Packet 3978: 7 -> 9 (AXI_WRITE)\n    inject_packet(7, 9, 64, "AXI_WRITE");\n    // Packet 3979: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 3980: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 827\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 827\n    // Packet 3981: 0 -> 12 (AXI_READ)\n    inject_packet(0, 12, 64, "AXI_READ");\n    // Packet 3982: 5 -> 0 (AXI_WRITE)\n    inject_packet(5, 0, 64, "AXI_WRITE");\n    // Packet 3983: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 3984: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 3985: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 3986: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 828\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 828\n    // Packet 3987: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 3988: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 3989: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 3990: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 3991: 9 -> 0 (AXI_WRITE)\n    inject_packet(9, 0, 64, "AXI_WRITE");\n    // Packet 3992: 11 -> 3 (AXI_READ)\n    inject_packet(11, 3, 64, "AXI_READ");\n    // Packet 3993: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 829\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 829\n    // Packet 3994: 5 -> 9 (AXI_READ)\n    inject_packet(5, 9, 64, "AXI_READ");\n    // Packet 3995: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 3996: 8 -> 14 (AXI_READ)\n    inject_packet(8, 14, 64, "AXI_READ");\n    // Packet 3997: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 831\n    repeat(2) @(posedge clk);\n    // Inject packets at cycle 831\n    // Packet 3998: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 3999: 1 -> 15 (AXI_WRITE)\n    inject_packet(1, 15, 64, "AXI_WRITE");\n    // Packet 4000: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 4001: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 4002: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 4003: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Packet 4004: 12 -> 0 (AXI_READ)\n    inject_packet(12, 0, 64, "AXI_READ");\n    // Wait until cycle 832\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 832\n    // Packet 4005: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Packet 4006: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 4007: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 4008: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 4009: 11 -> 2 (AXI_WRITE)\n    inject_packet(11, 2, 64, "AXI_WRITE");\n    // Wait until cycle 833\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 833\n    // Packet 4010: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 4011: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 4012: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 4013: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Wait until cycle 834\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 834\n    // Packet 4014: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 4015: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 4016: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 4017: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Wait until cycle 835\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 835\n    // Packet 4018: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 4019: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 4020: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 4021: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 4022: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 4023: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 4024: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Packet 4025: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 836\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 836\n    // Packet 4026: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 4027: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 4028: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Packet 4029: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 837\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 837\n    // Packet 4030: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 4031: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 4032: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 4033: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 4034: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 4035: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 838\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 838\n    // Packet 4036: 7 -> 2 (AXI_WRITE)\n    inject_packet(7, 2, 64, "AXI_WRITE");\n    // Wait until cycle 839\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 839\n    // Packet 4037: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 4038: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 4039: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Wait until cycle 840\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 840\n    // Packet 4040: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 4041: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 4042: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 4043: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 4044: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Wait until cycle 841\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 841\n    // Packet 4045: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 4046: 3 -> 14 (AXI_WRITE)\n    inject_packet(3, 14, 64, "AXI_WRITE");\n    // Packet 4047: 4 -> 3 (AXI_WRITE)\n    inject_packet(4, 3, 64, "AXI_WRITE");\n    // Packet 4048: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Wait until cycle 842\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 842\n    // Packet 4049: 1 -> 14 (AXI_READ)\n    inject_packet(1, 14, 64, "AXI_READ");\n    // Packet 4050: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 4051: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 4052: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Packet 4053: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Packet 4054: 11 -> 3 (AXI_WRITE)\n    inject_packet(11, 3, 64, "AXI_WRITE");\n    // Packet 4055: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Packet 4056: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 4057: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Packet 4058: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 843\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 843\n    // Packet 4059: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 4060: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 4061: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 4062: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 4063: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Packet 4064: 13 -> 5 (AXI_READ)\n    inject_packet(13, 5, 64, "AXI_READ");\n    // Packet 4065: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 844\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 844\n    // Packet 4066: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 4067: 6 -> 8 (AXI_WRITE)\n    inject_packet(6, 8, 64, "AXI_WRITE");\n    // Packet 4068: 7 -> 9 (AXI_READ)\n    inject_packet(7, 9, 64, "AXI_READ");\n    // Packet 4069: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 4070: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 845\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 845\n    // Packet 4071: 0 -> 4 (AXI_WRITE)\n    inject_packet(0, 4, 64, "AXI_WRITE");\n    // Packet 4072: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 4073: 8 -> 3 (AXI_WRITE)\n    inject_packet(8, 3, 64, "AXI_WRITE");\n    // Packet 4074: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 4075: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Packet 4076: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 846\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 846\n    // Packet 4077: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 4078: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 4079: 9 -> 13 (AXI_READ)\n    inject_packet(9, 13, 64, "AXI_READ");\n    // Packet 4080: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 4081: 11 -> 14 (AXI_READ)\n    inject_packet(11, 14, 64, "AXI_READ");\n    // Packet 4082: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Wait until cycle 847\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 847\n    // Packet 4083: 0 -> 11 (AXI_WRITE)\n    inject_packet(0, 11, 64, "AXI_WRITE");\n    // Packet 4084: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 4085: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Packet 4086: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 4087: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 848\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 848\n    // Packet 4088: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 4089: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 4090: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Packet 4091: 14 -> 0 (AXI_WRITE)\n    inject_packet(14, 0, 64, "AXI_WRITE");\n    // Wait until cycle 849\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 849\n    // Packet 4092: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 4093: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 4094: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Packet 4095: 15 -> 8 (AXI_READ)\n    inject_packet(15, 8, 64, "AXI_READ");\n    // Wait until cycle 850\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 850\n    // Packet 4096: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 4097: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 4098: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 4099: 9 -> 7 (AXI_READ)\n    inject_packet(9, 7, 64, "AXI_READ");\n    // Packet 4100: 14 -> 12 (AXI_READ)\n    inject_packet(14, 12, 64, "AXI_READ");\n    // Wait until cycle 851\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 851\n    // Packet 4101: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 4102: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 4103: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 4104: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 4105: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Wait until cycle 852\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 852\n    // Packet 4106: 2 -> 6 (AXI_READ)\n    inject_packet(2, 6, 64, "AXI_READ");\n    // Packet 4107: 4 -> 3 (AXI_READ)\n    inject_packet(4, 3, 64, "AXI_READ");\n    // Packet 4108: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 853\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 853\n    // Packet 4109: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 4110: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 4111: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 4112: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 854\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 854\n    // Packet 4113: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 4114: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 4115: 7 -> 9 (AXI_WRITE)\n    inject_packet(7, 9, 64, "AXI_WRITE");\n    // Packet 4116: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Wait until cycle 855\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 855\n    // Packet 4117: 1 -> 5 (AXI_WRITE)\n    inject_packet(1, 5, 64, "AXI_WRITE");\n    // Packet 4118: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 4119: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 4120: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Wait until cycle 856\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 856\n    // Packet 4121: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 4122: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 4123: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 4124: 6 -> 7 (AXI_READ)\n    inject_packet(6, 7, 64, "AXI_READ");\n    // Packet 4125: 9 -> 13 (AXI_WRITE)\n    inject_packet(9, 13, 64, "AXI_WRITE");\n    // Packet 4126: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 4127: 11 -> 6 (AXI_READ)\n    inject_packet(11, 6, 64, "AXI_READ");\n    // Packet 4128: 13 -> 0 (AXI_READ)\n    inject_packet(13, 0, 64, "AXI_READ");\n    // Packet 4129: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Wait until cycle 857\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 857\n    // Packet 4130: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 4131: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 4132: 8 -> 15 (AXI_WRITE)\n    inject_packet(8, 15, 64, "AXI_WRITE");\n    // Packet 4133: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 4134: 11 -> 5 (AXI_READ)\n    inject_packet(11, 5, 64, "AXI_READ");\n    // Packet 4135: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 858\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 858\n    // Packet 4136: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 4137: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 4138: 6 -> 7 (AXI_WRITE)\n    inject_packet(6, 7, 64, "AXI_WRITE");\n    // Packet 4139: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 4140: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 859\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 859\n    // Packet 4141: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 4142: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Packet 4143: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 4144: 9 -> 1 (AXI_WRITE)\n    inject_packet(9, 1, 64, "AXI_WRITE");\n    // Packet 4145: 10 -> 4 (AXI_WRITE)\n    inject_packet(10, 4, 64, "AXI_WRITE");\n    // Packet 4146: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Packet 4147: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 860\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 860\n    // Packet 4148: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 4149: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 4150: 7 -> 12 (AXI_READ)\n    inject_packet(7, 12, 64, "AXI_READ");\n    // Packet 4151: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 4152: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 4153: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Packet 4154: 15 -> 13 (AXI_WRITE)\n    inject_packet(15, 13, 64, "AXI_WRITE");\n    // Wait until cycle 861\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 861\n    // Packet 4155: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 4156: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 4157: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Packet 4158: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 862\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 862\n    // Packet 4159: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 4160: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 4161: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 4162: 12 -> 0 (AXI_WRITE)\n    inject_packet(12, 0, 64, "AXI_WRITE");\n    // Packet 4163: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Packet 4164: 15 -> 2 (AXI_WRITE)\n    inject_packet(15, 2, 64, "AXI_WRITE");\n    // Wait until cycle 863\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 863\n    // Packet 4165: 1 -> 3 (AXI_READ)\n    inject_packet(1, 3, 64, "AXI_READ");\n    // Packet 4166: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 4167: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 4168: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 4169: 9 -> 13 (AXI_READ)\n    inject_packet(9, 13, 64, "AXI_READ");\n    // Packet 4170: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 4171: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 4172: 13 -> 2 (AXI_WRITE)\n    inject_packet(13, 2, 64, "AXI_WRITE");\n    // Wait until cycle 864\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 864\n    // Packet 4173: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 4174: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 4175: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Packet 4176: 8 -> 15 (AXI_READ)\n    inject_packet(8, 15, 64, "AXI_READ");\n    // Packet 4177: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 865\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 865\n    // Packet 4178: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 4179: 1 -> 8 (AXI_WRITE)\n    inject_packet(1, 8, 64, "AXI_WRITE");\n    // Packet 4180: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 4181: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Packet 4182: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 866\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 866\n    // Packet 4183: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 4184: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 4185: 8 -> 1 (AXI_READ)\n    inject_packet(8, 1, 64, "AXI_READ");\n    // Packet 4186: 14 -> 9 (AXI_READ)\n    inject_packet(14, 9, 64, "AXI_READ");\n    // Wait until cycle 867\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 867\n    // Packet 4187: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 4188: 4 -> 1 (AXI_READ)\n    inject_packet(4, 1, 64, "AXI_READ");\n    // Packet 4189: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 4190: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 4191: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 4192: 9 -> 11 (AXI_READ)\n    inject_packet(9, 11, 64, "AXI_READ");\n    // Packet 4193: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 4194: 15 -> 7 (AXI_READ)\n    inject_packet(15, 7, 64, "AXI_READ");\n    // Wait until cycle 868\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 868\n    // Packet 4195: 3 -> 1 (AXI_READ)\n    inject_packet(3, 1, 64, "AXI_READ");\n    // Packet 4196: 5 -> 13 (AXI_WRITE)\n    inject_packet(5, 13, 64, "AXI_WRITE");\n    // Packet 4197: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 4198: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 869\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 869\n    // Packet 4199: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 4200: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 4201: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 4202: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Wait until cycle 870\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 870\n    // Packet 4203: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 4204: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 4205: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Packet 4206: 14 -> 13 (AXI_WRITE)\n    inject_packet(14, 13, 64, "AXI_WRITE");\n    // Packet 4207: 15 -> 1 (AXI_READ)\n    inject_packet(15, 1, 64, "AXI_READ");\n    // Wait until cycle 871\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 871\n    // Packet 4208: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Packet 4209: 11 -> 2 (AXI_READ)\n    inject_packet(11, 2, 64, "AXI_READ");\n    // Packet 4210: 12 -> 4 (AXI_READ)\n    inject_packet(12, 4, 64, "AXI_READ");\n    // Packet 4211: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 872\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 872\n    // Packet 4212: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 4213: 6 -> 14 (AXI_WRITE)\n    inject_packet(6, 14, 64, "AXI_WRITE");\n    // Packet 4214: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 4215: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 4216: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 4217: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Packet 4218: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 873\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 873\n    // Packet 4219: 1 -> 3 (AXI_WRITE)\n    inject_packet(1, 3, 64, "AXI_WRITE");\n    // Packet 4220: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 4221: 5 -> 0 (AXI_WRITE)\n    inject_packet(5, 0, 64, "AXI_WRITE");\n    // Packet 4222: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 4223: 10 -> 1 (AXI_WRITE)\n    inject_packet(10, 1, 64, "AXI_WRITE");\n    // Packet 4224: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 4225: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Packet 4226: 15 -> 9 (AXI_WRITE)\n    inject_packet(15, 9, 64, "AXI_WRITE");\n    // Wait until cycle 874\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 874\n    // Packet 4227: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 4228: 1 -> 2 (AXI_WRITE)\n    inject_packet(1, 2, 64, "AXI_WRITE");\n    // Packet 4229: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 4230: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 4231: 9 -> 1 (AXI_WRITE)\n    inject_packet(9, 1, 64, "AXI_WRITE");\n    // Packet 4232: 10 -> 3 (AXI_READ)\n    inject_packet(10, 3, 64, "AXI_READ");\n    // Packet 4233: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Packet 4234: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Wait until cycle 875\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 875\n    // Packet 4235: 10 -> 0 (AXI_WRITE)\n    inject_packet(10, 0, 64, "AXI_WRITE");\n    // Packet 4236: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 876\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 876\n    // Packet 4237: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 4238: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 4239: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 4240: 7 -> 4 (AXI_READ)\n    inject_packet(7, 4, 64, "AXI_READ");\n    // Packet 4241: 9 -> 4 (AXI_WRITE)\n    inject_packet(9, 4, 64, "AXI_WRITE");\n    // Packet 4242: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Wait until cycle 877\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 877\n    // Packet 4243: 0 -> 6 (AXI_WRITE)\n    inject_packet(0, 6, 64, "AXI_WRITE");\n    // Packet 4244: 3 -> 14 (AXI_READ)\n    inject_packet(3, 14, 64, "AXI_READ");\n    // Packet 4245: 6 -> 8 (AXI_READ)\n    inject_packet(6, 8, 64, "AXI_READ");\n    // Packet 4246: 7 -> 6 (AXI_WRITE)\n    inject_packet(7, 6, 64, "AXI_WRITE");\n    // Packet 4247: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Packet 4248: 10 -> 14 (AXI_WRITE)\n    inject_packet(10, 14, 64, "AXI_WRITE");\n    // Packet 4249: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Wait until cycle 878\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 878\n    // Packet 4250: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 4251: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 4252: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 4253: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 4254: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 4255: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Wait until cycle 879\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 879\n    // Packet 4256: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 4257: 1 -> 15 (AXI_WRITE)\n    inject_packet(1, 15, 64, "AXI_WRITE");\n    // Packet 4258: 8 -> 12 (AXI_READ)\n    inject_packet(8, 12, 64, "AXI_READ");\n    // Packet 4259: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Wait until cycle 880\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 880\n    // Packet 4260: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 4261: 6 -> 3 (AXI_WRITE)\n    inject_packet(6, 3, 64, "AXI_WRITE");\n    // Packet 4262: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 4263: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Packet 4264: 11 -> 6 (AXI_READ)\n    inject_packet(11, 6, 64, "AXI_READ");\n    // Packet 4265: 12 -> 6 (AXI_WRITE)\n    inject_packet(12, 6, 64, "AXI_WRITE");\n    // Packet 4266: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 881\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 881\n    // Packet 4267: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 4268: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 4269: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 882\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 882\n    // Packet 4270: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 4271: 3 -> 11 (AXI_READ)\n    inject_packet(3, 11, 64, "AXI_READ");\n    // Packet 4272: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 883\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 883\n    // Packet 4273: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 4274: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 4275: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 4276: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Packet 4277: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 4278: 14 -> 13 (AXI_READ)\n    inject_packet(14, 13, 64, "AXI_READ");\n    // Wait until cycle 884\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 884\n    // Packet 4279: 2 -> 1 (AXI_READ)\n    inject_packet(2, 1, 64, "AXI_READ");\n    // Packet 4280: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 4281: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 4282: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Packet 4283: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Packet 4284: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 885\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 885\n    // Packet 4285: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 4286: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 4287: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 4288: 10 -> 5 (AXI_WRITE)\n    inject_packet(10, 5, 64, "AXI_WRITE");\n    // Packet 4289: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Wait until cycle 886\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 886\n    // Packet 4290: 0 -> 1 (AXI_READ)\n    inject_packet(0, 1, 64, "AXI_READ");\n    // Packet 4291: 4 -> 12 (AXI_READ)\n    inject_packet(4, 12, 64, "AXI_READ");\n    // Wait until cycle 887\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 887\n    // Packet 4292: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 4293: 6 -> 14 (AXI_READ)\n    inject_packet(6, 14, 64, "AXI_READ");\n    // Packet 4294: 8 -> 7 (AXI_READ)\n    inject_packet(8, 7, 64, "AXI_READ");\n    // Packet 4295: 9 -> 0 (AXI_READ)\n    inject_packet(9, 0, 64, "AXI_READ");\n    // Packet 4296: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Packet 4297: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Wait until cycle 888\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 888\n    // Packet 4298: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 4299: 1 -> 3 (AXI_WRITE)\n    inject_packet(1, 3, 64, "AXI_WRITE");\n    // Packet 4300: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 4301: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Packet 4302: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 889\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 889\n    // Packet 4303: 1 -> 10 (AXI_WRITE)\n    inject_packet(1, 10, 64, "AXI_WRITE");\n    // Packet 4304: 3 -> 8 (AXI_WRITE)\n    inject_packet(3, 8, 64, "AXI_WRITE");\n    // Packet 4305: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 4306: 7 -> 1 (AXI_WRITE)\n    inject_packet(7, 1, 64, "AXI_WRITE");\n    // Packet 4307: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 4308: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Wait until cycle 890\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 890\n    // Packet 4309: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 4310: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 4311: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 4312: 10 -> 9 (AXI_READ)\n    inject_packet(10, 9, 64, "AXI_READ");\n    // Packet 4313: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Packet 4314: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 891\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 891\n    // Packet 4315: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 4316: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 4317: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 4318: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 4319: 12 -> 13 (AXI_READ)\n    inject_packet(12, 13, 64, "AXI_READ");\n    // Wait until cycle 892\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 892\n    // Packet 4320: 1 -> 0 (AXI_READ)\n    inject_packet(1, 0, 64, "AXI_READ");\n    // Packet 4321: 4 -> 15 (AXI_READ)\n    inject_packet(4, 15, 64, "AXI_READ");\n    // Packet 4322: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 4323: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 4324: 10 -> 3 (AXI_READ)\n    inject_packet(10, 3, 64, "AXI_READ");\n    // Packet 4325: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Wait until cycle 893\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 893\n    // Packet 4326: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 4327: 8 -> 0 (AXI_WRITE)\n    inject_packet(8, 0, 64, "AXI_WRITE");\n    // Packet 4328: 9 -> 8 (AXI_WRITE)\n    inject_packet(9, 8, 64, "AXI_WRITE");\n    // Packet 4329: 10 -> 6 (AXI_READ)\n    inject_packet(10, 6, 64, "AXI_READ");\n    // Packet 4330: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Packet 4331: 12 -> 7 (AXI_WRITE)\n    inject_packet(12, 7, 64, "AXI_WRITE");\n    // Packet 4332: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Wait until cycle 894\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 894\n    // Packet 4333: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 4334: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 4335: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 4336: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 4337: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 4338: 15 -> 9 (AXI_READ)\n    inject_packet(15, 9, 64, "AXI_READ");\n    // Wait until cycle 895\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 895\n    // Packet 4339: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 4340: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 4341: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 4342: 5 -> 0 (AXI_WRITE)\n    inject_packet(5, 0, 64, "AXI_WRITE");\n    // Packet 4343: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 4344: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Packet 4345: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Packet 4346: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 896\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 896\n    // Packet 4347: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 4348: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 4349: 9 -> 0 (AXI_WRITE)\n    inject_packet(9, 0, 64, "AXI_WRITE");\n    // Packet 4350: 12 -> 8 (AXI_READ)\n    inject_packet(12, 8, 64, "AXI_READ");\n    // Packet 4351: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Packet 4352: 14 -> 15 (AXI_WRITE)\n    inject_packet(14, 15, 64, "AXI_WRITE");\n    // Wait until cycle 897\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 897\n    // Packet 4353: 2 -> 5 (AXI_WRITE)\n    inject_packet(2, 5, 64, "AXI_WRITE");\n    // Packet 4354: 3 -> 10 (AXI_READ)\n    inject_packet(3, 10, 64, "AXI_READ");\n    // Packet 4355: 7 -> 0 (AXI_READ)\n    inject_packet(7, 0, 64, "AXI_READ");\n    // Packet 4356: 11 -> 9 (AXI_WRITE)\n    inject_packet(11, 9, 64, "AXI_WRITE");\n    // Wait until cycle 898\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 898\n    // Packet 4357: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 4358: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Wait until cycle 899\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 899\n    // Packet 4359: 0 -> 1 (AXI_WRITE)\n    inject_packet(0, 1, 64, "AXI_WRITE");\n    // Packet 4360: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 4361: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 4362: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Wait until cycle 900\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 900\n    // Packet 4363: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 4364: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 4365: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Packet 4366: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 4367: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 901\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 901\n    // Packet 4368: 9 -> 12 (AXI_READ)\n    inject_packet(9, 12, 64, "AXI_READ");\n    // Packet 4369: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 4370: 12 -> 5 (AXI_WRITE)\n    inject_packet(12, 5, 64, "AXI_WRITE");\n    // Packet 4371: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 4372: 15 -> 12 (AXI_WRITE)\n    inject_packet(15, 12, 64, "AXI_WRITE");\n    // Wait until cycle 902\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 902\n    // Packet 4373: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 4374: 6 -> 12 (AXI_WRITE)\n    inject_packet(6, 12, 64, "AXI_WRITE");\n    // Packet 4375: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 4376: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 4377: 11 -> 4 (AXI_READ)\n    inject_packet(11, 4, 64, "AXI_READ");\n    // Wait until cycle 903\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 903\n    // Packet 4378: 5 -> 15 (AXI_READ)\n    inject_packet(5, 15, 64, "AXI_READ");\n    // Packet 4379: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 4380: 10 -> 12 (AXI_READ)\n    inject_packet(10, 12, 64, "AXI_READ");\n    // Packet 4381: 11 -> 5 (AXI_WRITE)\n    inject_packet(11, 5, 64, "AXI_WRITE");\n    // Packet 4382: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Wait until cycle 904\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 904\n    // Packet 4383: 0 -> 7 (AXI_WRITE)\n    inject_packet(0, 7, 64, "AXI_WRITE");\n    // Packet 4384: 1 -> 12 (AXI_WRITE)\n    inject_packet(1, 12, 64, "AXI_WRITE");\n    // Packet 4385: 2 -> 15 (AXI_WRITE)\n    inject_packet(2, 15, 64, "AXI_WRITE");\n    // Packet 4386: 3 -> 7 (AXI_READ)\n    inject_packet(3, 7, 64, "AXI_READ");\n    // Packet 4387: 8 -> 15 (AXI_READ)\n    inject_packet(8, 15, 64, "AXI_READ");\n    // Packet 4388: 11 -> 0 (AXI_READ)\n    inject_packet(11, 0, 64, "AXI_READ");\n    // Wait until cycle 905\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 905\n    // Packet 4389: 3 -> 2 (AXI_READ)\n    inject_packet(3, 2, 64, "AXI_READ");\n    // Packet 4390: 12 -> 3 (AXI_READ)\n    inject_packet(12, 3, 64, "AXI_READ");\n    // Packet 4391: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Wait until cycle 906\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 906\n    // Packet 4392: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 4393: 5 -> 11 (AXI_READ)\n    inject_packet(5, 11, 64, "AXI_READ");\n    // Packet 4394: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 4395: 7 -> 8 (AXI_READ)\n    inject_packet(7, 8, 64, "AXI_READ");\n    // Packet 4396: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 4397: 11 -> 7 (AXI_WRITE)\n    inject_packet(11, 7, 64, "AXI_WRITE");\n    // Packet 4398: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Wait until cycle 907\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 907\n    // Packet 4399: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 4400: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 4401: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 4402: 12 -> 6 (AXI_READ)\n    inject_packet(12, 6, 64, "AXI_READ");\n    // Packet 4403: 13 -> 11 (AXI_WRITE)\n    inject_packet(13, 11, 64, "AXI_WRITE");\n    // Wait until cycle 908\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 908\n    // Packet 4404: 1 -> 7 (AXI_READ)\n    inject_packet(1, 7, 64, "AXI_READ");\n    // Packet 4405: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 4406: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 4407: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 4408: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 4409: 11 -> 0 (AXI_READ)\n    inject_packet(11, 0, 64, "AXI_READ");\n    // Packet 4410: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Packet 4411: 15 -> 0 (AXI_READ)\n    inject_packet(15, 0, 64, "AXI_READ");\n    // Wait until cycle 909\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 909\n    // Packet 4412: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 4413: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 4414: 5 -> 2 (AXI_READ)\n    inject_packet(5, 2, 64, "AXI_READ");\n    // Packet 4415: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Wait until cycle 910\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 910\n    // Packet 4416: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 4417: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 4418: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 4419: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 4420: 12 -> 4 (AXI_WRITE)\n    inject_packet(12, 4, 64, "AXI_WRITE");\n    // Packet 4421: 13 -> 1 (AXI_READ)\n    inject_packet(13, 1, 64, "AXI_READ");\n    // Wait until cycle 911\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 911\n    // Packet 4422: 0 -> 9 (AXI_WRITE)\n    inject_packet(0, 9, 64, "AXI_WRITE");\n    // Packet 4423: 3 -> 15 (AXI_WRITE)\n    inject_packet(3, 15, 64, "AXI_WRITE");\n    // Packet 4424: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 4425: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 4426: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Packet 4427: 14 -> 6 (AXI_READ)\n    inject_packet(14, 6, 64, "AXI_READ");\n    // Wait until cycle 912\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 912\n    // Packet 4428: 2 -> 14 (AXI_READ)\n    inject_packet(2, 14, 64, "AXI_READ");\n    // Packet 4429: 6 -> 5 (AXI_READ)\n    inject_packet(6, 5, 64, "AXI_READ");\n    // Packet 4430: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Packet 4431: 10 -> 3 (AXI_READ)\n    inject_packet(10, 3, 64, "AXI_READ");\n    // Packet 4432: 14 -> 8 (AXI_WRITE)\n    inject_packet(14, 8, 64, "AXI_WRITE");\n    // Wait until cycle 913\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 913\n    // Packet 4433: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 4434: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 4435: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Packet 4436: 8 -> 13 (AXI_WRITE)\n    inject_packet(8, 13, 64, "AXI_WRITE");\n    // Packet 4437: 12 -> 11 (AXI_WRITE)\n    inject_packet(12, 11, 64, "AXI_WRITE");\n    // Packet 4438: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 914\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 914\n    // Packet 4439: 9 -> 3 (AXI_READ)\n    inject_packet(9, 3, 64, "AXI_READ");\n    // Wait until cycle 915\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 915\n    // Packet 4440: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 4441: 12 -> 2 (AXI_READ)\n    inject_packet(12, 2, 64, "AXI_READ");\n    // Packet 4442: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Packet 4443: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 916\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 916\n    // Packet 4444: 4 -> 10 (AXI_WRITE)\n    inject_packet(4, 10, 64, "AXI_WRITE");\n    // Packet 4445: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Wait until cycle 917\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 917\n    // Packet 4446: 0 -> 3 (AXI_WRITE)\n    inject_packet(0, 3, 64, "AXI_WRITE");\n    // Packet 4447: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 4448: 3 -> 9 (AXI_WRITE)\n    inject_packet(3, 9, 64, "AXI_WRITE");\n    // Packet 4449: 5 -> 3 (AXI_READ)\n    inject_packet(5, 3, 64, "AXI_READ");\n    // Packet 4450: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 4451: 8 -> 6 (AXI_READ)\n    inject_packet(8, 6, 64, "AXI_READ");\n    // Packet 4452: 9 -> 13 (AXI_READ)\n    inject_packet(9, 13, 64, "AXI_READ");\n    // Packet 4453: 11 -> 3 (AXI_WRITE)\n    inject_packet(11, 3, 64, "AXI_WRITE");\n    // Packet 4454: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Packet 4455: 15 -> 10 (AXI_WRITE)\n    inject_packet(15, 10, 64, "AXI_WRITE");\n    // Wait until cycle 918\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 918\n    // Packet 4456: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 4457: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 4458: 10 -> 3 (AXI_READ)\n    inject_packet(10, 3, 64, "AXI_READ");\n    // Packet 4459: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 4460: 14 -> 2 (AXI_READ)\n    inject_packet(14, 2, 64, "AXI_READ");\n    // Wait until cycle 919\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 919\n    // Packet 4461: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 4462: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 4463: 15 -> 5 (AXI_READ)\n    inject_packet(15, 5, 64, "AXI_READ");\n    // Wait until cycle 920\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 920\n    // Packet 4464: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 4465: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 4466: 7 -> 8 (AXI_WRITE)\n    inject_packet(7, 8, 64, "AXI_WRITE");\n    // Packet 4467: 9 -> 7 (AXI_WRITE)\n    inject_packet(9, 7, 64, "AXI_WRITE");\n    // Packet 4468: 10 -> 11 (AXI_WRITE)\n    inject_packet(10, 11, 64, "AXI_WRITE");\n    // Wait until cycle 921\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 921\n    // Packet 4469: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 4470: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 4471: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 4472: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Wait until cycle 922\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 922\n    // Packet 4473: 2 -> 15 (AXI_READ)\n    inject_packet(2, 15, 64, "AXI_READ");\n    // Packet 4474: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 4475: 10 -> 15 (AXI_WRITE)\n    inject_packet(10, 15, 64, "AXI_WRITE");\n    // Packet 4476: 11 -> 12 (AXI_WRITE)\n    inject_packet(11, 12, 64, "AXI_WRITE");\n    // Packet 4477: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 4478: 14 -> 6 (AXI_WRITE)\n    inject_packet(14, 6, 64, "AXI_WRITE");\n    // Packet 4479: 15 -> 2 (AXI_READ)\n    inject_packet(15, 2, 64, "AXI_READ");\n    // Wait until cycle 923\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 923\n    // Packet 4480: 2 -> 7 (AXI_READ)\n    inject_packet(2, 7, 64, "AXI_READ");\n    // Packet 4481: 3 -> 2 (AXI_READ)\n    inject_packet(3, 2, 64, "AXI_READ");\n    // Packet 4482: 7 -> 15 (AXI_WRITE)\n    inject_packet(7, 15, 64, "AXI_WRITE");\n    // Packet 4483: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Packet 4484: 10 -> 7 (AXI_WRITE)\n    inject_packet(10, 7, 64, "AXI_WRITE");\n    // Packet 4485: 14 -> 3 (AXI_WRITE)\n    inject_packet(14, 3, 64, "AXI_WRITE");\n    // Wait until cycle 924\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 924\n    // Packet 4486: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 4487: 6 -> 9 (AXI_READ)\n    inject_packet(6, 9, 64, "AXI_READ");\n    // Packet 4488: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 4489: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 4490: 10 -> 8 (AXI_READ)\n    inject_packet(10, 8, 64, "AXI_READ");\n    // Packet 4491: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 4492: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 925\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 925\n    // Packet 4493: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 4494: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Wait until cycle 926\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 926\n    // Packet 4495: 0 -> 13 (AXI_READ)\n    inject_packet(0, 13, 64, "AXI_READ");\n    // Packet 4496: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 4497: 3 -> 1 (AXI_WRITE)\n    inject_packet(3, 1, 64, "AXI_WRITE");\n    // Packet 4498: 5 -> 7 (AXI_WRITE)\n    inject_packet(5, 7, 64, "AXI_WRITE");\n    // Wait until cycle 927\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 927\n    // Packet 4499: 4 -> 8 (AXI_WRITE)\n    inject_packet(4, 8, 64, "AXI_WRITE");\n    // Packet 4500: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 4501: 12 -> 0 (AXI_WRITE)\n    inject_packet(12, 0, 64, "AXI_WRITE");\n    // Packet 4502: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Packet 4503: 14 -> 1 (AXI_READ)\n    inject_packet(14, 1, 64, "AXI_READ");\n    // Packet 4504: 15 -> 4 (AXI_WRITE)\n    inject_packet(15, 4, 64, "AXI_WRITE");\n    // Wait until cycle 928\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 928\n    // Packet 4505: 0 -> 13 (AXI_WRITE)\n    inject_packet(0, 13, 64, "AXI_WRITE");\n    // Packet 4506: 2 -> 13 (AXI_READ)\n    inject_packet(2, 13, 64, "AXI_READ");\n    // Packet 4507: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 4508: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 4509: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Packet 4510: 14 -> 15 (AXI_READ)\n    inject_packet(14, 15, 64, "AXI_READ");\n    // Wait until cycle 929\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 929\n    // Packet 4511: 1 -> 13 (AXI_WRITE)\n    inject_packet(1, 13, 64, "AXI_WRITE");\n    // Packet 4512: 5 -> 10 (AXI_WRITE)\n    inject_packet(5, 10, 64, "AXI_WRITE");\n    // Packet 4513: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 4514: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Wait until cycle 930\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 930\n    // Packet 4515: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 4516: 3 -> 6 (AXI_WRITE)\n    inject_packet(3, 6, 64, "AXI_WRITE");\n    // Packet 4517: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Packet 4518: 14 -> 5 (AXI_WRITE)\n    inject_packet(14, 5, 64, "AXI_WRITE");\n    // Wait until cycle 931\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 931\n    // Packet 4519: 7 -> 6 (AXI_READ)\n    inject_packet(7, 6, 64, "AXI_READ");\n    // Packet 4520: 8 -> 10 (AXI_WRITE)\n    inject_packet(8, 10, 64, "AXI_WRITE");\n    // Packet 4521: 9 -> 11 (AXI_READ)\n    inject_packet(9, 11, 64, "AXI_READ");\n    // Packet 4522: 15 -> 8 (AXI_WRITE)\n    inject_packet(15, 8, 64, "AXI_WRITE");\n    // Wait until cycle 932\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 932\n    // Packet 4523: 4 -> 3 (AXI_READ)\n    inject_packet(4, 3, 64, "AXI_READ");\n    // Packet 4524: 8 -> 6 (AXI_WRITE)\n    inject_packet(8, 6, 64, "AXI_WRITE");\n    // Packet 4525: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Wait until cycle 933\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 933\n    // Packet 4526: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 4527: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 4528: 10 -> 11 (AXI_READ)\n    inject_packet(10, 11, 64, "AXI_READ");\n    // Packet 4529: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Packet 4530: 12 -> 10 (AXI_WRITE)\n    inject_packet(12, 10, 64, "AXI_WRITE");\n    // Wait until cycle 934\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 934\n    // Packet 4531: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 4532: 2 -> 9 (AXI_READ)\n    inject_packet(2, 9, 64, "AXI_READ");\n    // Packet 4533: 3 -> 8 (AXI_READ)\n    inject_packet(3, 8, 64, "AXI_READ");\n    // Packet 4534: 6 -> 10 (AXI_READ)\n    inject_packet(6, 10, 64, "AXI_READ");\n    // Wait until cycle 935\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 935\n    // Packet 4535: 1 -> 3 (AXI_WRITE)\n    inject_packet(1, 3, 64, "AXI_WRITE");\n    // Packet 4536: 10 -> 7 (AXI_READ)\n    inject_packet(10, 7, 64, "AXI_READ");\n    // Packet 4537: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n    // Wait until cycle 936\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 936\n    // Packet 4538: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 4539: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 4540: 4 -> 13 (AXI_WRITE)\n    inject_packet(4, 13, 64, "AXI_WRITE");\n    // Packet 4541: 5 -> 15 (AXI_WRITE)\n    inject_packet(5, 15, 64, "AXI_WRITE");\n    // Packet 4542: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 4543: 13 -> 8 (AXI_READ)\n    inject_packet(13, 8, 64, "AXI_READ");\n    // Wait until cycle 937\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 937\n    // Packet 4544: 2 -> 8 (AXI_READ)\n    inject_packet(2, 8, 64, "AXI_READ");\n    // Packet 4545: 4 -> 10 (AXI_READ)\n    inject_packet(4, 10, 64, "AXI_READ");\n    // Wait until cycle 938\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 938\n    // Packet 4546: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 4547: 6 -> 10 (AXI_WRITE)\n    inject_packet(6, 10, 64, "AXI_WRITE");\n    // Packet 4548: 8 -> 15 (AXI_READ)\n    inject_packet(8, 15, 64, "AXI_READ");\n    // Packet 4549: 11 -> 15 (AXI_READ)\n    inject_packet(11, 15, 64, "AXI_READ");\n    // Packet 4550: 12 -> 9 (AXI_WRITE)\n    inject_packet(12, 9, 64, "AXI_WRITE");\n    // Packet 4551: 15 -> 12 (AXI_READ)\n    inject_packet(15, 12, 64, "AXI_READ");\n    // Wait until cycle 939\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 939\n    // Packet 4552: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 4553: 2 -> 7 (AXI_WRITE)\n    inject_packet(2, 7, 64, "AXI_WRITE");\n    // Packet 4554: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 4555: 8 -> 13 (AXI_READ)\n    inject_packet(8, 13, 64, "AXI_READ");\n    // Packet 4556: 10 -> 8 (AXI_READ)\n    inject_packet(10, 8, 64, "AXI_READ");\n    // Packet 4557: 11 -> 15 (AXI_WRITE)\n    inject_packet(11, 15, 64, "AXI_WRITE");\n    // Packet 4558: 15 -> 11 (AXI_WRITE)\n    inject_packet(15, 11, 64, "AXI_WRITE");\n    // Wait until cycle 940\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 940\n    // Packet 4559: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 4560: 7 -> 5 (AXI_WRITE)\n    inject_packet(7, 5, 64, "AXI_WRITE");\n    // Packet 4561: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 4562: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Packet 4563: 13 -> 5 (AXI_WRITE)\n    inject_packet(13, 5, 64, "AXI_WRITE");\n    // Wait until cycle 941\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 941\n    // Packet 4564: 11 -> 0 (AXI_WRITE)\n    inject_packet(11, 0, 64, "AXI_WRITE");\n    // Packet 4565: 14 -> 1 (AXI_WRITE)\n    inject_packet(14, 1, 64, "AXI_WRITE");\n    // Packet 4566: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 942\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 942\n    // Packet 4567: 8 -> 9 (AXI_WRITE)\n    inject_packet(8, 9, 64, "AXI_WRITE");\n    // Packet 4568: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Wait until cycle 943\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 943\n    // Packet 4569: 4 -> 11 (AXI_WRITE)\n    inject_packet(4, 11, 64, "AXI_WRITE");\n    // Packet 4570: 9 -> 7 (AXI_WRITE)\n    inject_packet(9, 7, 64, "AXI_WRITE");\n    // Packet 4571: 10 -> 13 (AXI_READ)\n    inject_packet(10, 13, 64, "AXI_READ");\n    // Wait until cycle 944\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 944\n    // Packet 4572: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 4573: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 4574: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 4575: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 4576: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 945\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 945\n    // Packet 4577: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 4578: 5 -> 4 (AXI_READ)\n    inject_packet(5, 4, 64, "AXI_READ");\n    // Packet 4579: 11 -> 3 (AXI_WRITE)\n    inject_packet(11, 3, 64, "AXI_WRITE");\n    // Packet 4580: 13 -> 7 (AXI_READ)\n    inject_packet(13, 7, 64, "AXI_READ");\n    // Packet 4581: 14 -> 12 (AXI_WRITE)\n    inject_packet(14, 12, 64, "AXI_WRITE");\n    // Wait until cycle 946\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 946\n    // Packet 4582: 6 -> 1 (AXI_WRITE)\n    inject_packet(6, 1, 64, "AXI_WRITE");\n    // Packet 4583: 7 -> 15 (AXI_READ)\n    inject_packet(7, 15, 64, "AXI_READ");\n    // Packet 4584: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Wait until cycle 947\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 947\n    // Packet 4585: 3 -> 13 (AXI_WRITE)\n    inject_packet(3, 13, 64, "AXI_WRITE");\n    // Packet 4586: 9 -> 8 (AXI_READ)\n    inject_packet(9, 8, 64, "AXI_READ");\n    // Packet 4587: 12 -> 11 (AXI_READ)\n    inject_packet(12, 11, 64, "AXI_READ");\n    // Packet 4588: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 948\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 948\n    // Packet 4589: 4 -> 2 (AXI_WRITE)\n    inject_packet(4, 2, 64, "AXI_WRITE");\n    // Packet 4590: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 949\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 949\n    // Packet 4591: 0 -> 12 (AXI_WRITE)\n    inject_packet(0, 12, 64, "AXI_WRITE");\n    // Packet 4592: 4 -> 6 (AXI_WRITE)\n    inject_packet(4, 6, 64, "AXI_WRITE");\n    // Packet 4593: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 4594: 7 -> 14 (AXI_READ)\n    inject_packet(7, 14, 64, "AXI_READ");\n    // Packet 4595: 8 -> 12 (AXI_READ)\n    inject_packet(8, 12, 64, "AXI_READ");\n    // Packet 4596: 9 -> 10 (AXI_READ)\n    inject_packet(9, 10, 64, "AXI_READ");\n    // Packet 4597: 10 -> 3 (AXI_WRITE)\n    inject_packet(10, 3, 64, "AXI_WRITE");\n    // Wait until cycle 950\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 950\n    // Packet 4598: 0 -> 8 (AXI_WRITE)\n    inject_packet(0, 8, 64, "AXI_WRITE");\n    // Packet 4599: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 4600: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 4601: 6 -> 13 (AXI_WRITE)\n    inject_packet(6, 13, 64, "AXI_WRITE");\n    // Packet 4602: 7 -> 4 (AXI_WRITE)\n    inject_packet(7, 4, 64, "AXI_WRITE");\n    // Packet 4603: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Packet 4604: 14 -> 12 (AXI_READ)\n    inject_packet(14, 12, 64, "AXI_READ");\n    // Wait until cycle 951\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 951\n    // Packet 4605: 0 -> 10 (AXI_WRITE)\n    inject_packet(0, 10, 64, "AXI_WRITE");\n    // Packet 4606: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Packet 4607: 13 -> 15 (AXI_WRITE)\n    inject_packet(13, 15, 64, "AXI_WRITE");\n    // Packet 4608: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Wait until cycle 952\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 952\n    // Packet 4609: 4 -> 5 (AXI_WRITE)\n    inject_packet(4, 5, 64, "AXI_WRITE");\n    // Packet 4610: 7 -> 9 (AXI_READ)\n    inject_packet(7, 9, 64, "AXI_READ");\n    // Packet 4611: 12 -> 15 (AXI_WRITE)\n    inject_packet(12, 15, 64, "AXI_WRITE");\n    // Packet 4612: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Wait until cycle 953\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 953\n    // Packet 4613: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 4614: 2 -> 12 (AXI_WRITE)\n    inject_packet(2, 12, 64, "AXI_WRITE");\n    // Packet 4615: 6 -> 2 (AXI_READ)\n    inject_packet(6, 2, 64, "AXI_READ");\n    // Packet 4616: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 4617: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 4618: 12 -> 8 (AXI_WRITE)\n    inject_packet(12, 8, 64, "AXI_WRITE");\n    // Packet 4619: 14 -> 11 (AXI_WRITE)\n    inject_packet(14, 11, 64, "AXI_WRITE");\n    // Wait until cycle 954\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 954\n    // Packet 4620: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 4621: 3 -> 7 (AXI_WRITE)\n    inject_packet(3, 7, 64, "AXI_WRITE");\n    // Packet 4622: 5 -> 1 (AXI_READ)\n    inject_packet(5, 1, 64, "AXI_READ");\n    // Packet 4623: 9 -> 10 (AXI_WRITE)\n    inject_packet(9, 10, 64, "AXI_WRITE");\n    // Packet 4624: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 955\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 955\n    // Packet 4625: 0 -> 7 (AXI_READ)\n    inject_packet(0, 7, 64, "AXI_READ");\n    // Packet 4626: 1 -> 13 (AXI_READ)\n    inject_packet(1, 13, 64, "AXI_READ");\n    // Packet 4627: 3 -> 12 (AXI_READ)\n    inject_packet(3, 12, 64, "AXI_READ");\n    // Packet 4628: 4 -> 0 (AXI_READ)\n    inject_packet(4, 0, 64, "AXI_READ");\n    // Packet 4629: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 4630: 12 -> 5 (AXI_READ)\n    inject_packet(12, 5, 64, "AXI_READ");\n    // Packet 4631: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Packet 4632: 14 -> 12 (AXI_READ)\n    inject_packet(14, 12, 64, "AXI_READ");\n    // Packet 4633: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 956\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 956\n    // Packet 4634: 0 -> 6 (AXI_READ)\n    inject_packet(0, 6, 64, "AXI_READ");\n    // Packet 4635: 1 -> 12 (AXI_READ)\n    inject_packet(1, 12, 64, "AXI_READ");\n    // Packet 4636: 2 -> 14 (AXI_WRITE)\n    inject_packet(2, 14, 64, "AXI_WRITE");\n    // Packet 4637: 4 -> 14 (AXI_READ)\n    inject_packet(4, 14, 64, "AXI_READ");\n    // Packet 4638: 5 -> 14 (AXI_READ)\n    inject_packet(5, 14, 64, "AXI_READ");\n    // Packet 4639: 6 -> 0 (AXI_WRITE)\n    inject_packet(6, 0, 64, "AXI_WRITE");\n    // Packet 4640: 7 -> 10 (AXI_READ)\n    inject_packet(7, 10, 64, "AXI_READ");\n    // Packet 4641: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 4642: 10 -> 0 (AXI_READ)\n    inject_packet(10, 0, 64, "AXI_READ");\n    // Packet 4643: 15 -> 3 (AXI_WRITE)\n    inject_packet(15, 3, 64, "AXI_WRITE");\n    // Wait until cycle 957\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 957\n    // Packet 4644: 1 -> 10 (AXI_READ)\n    inject_packet(1, 10, 64, "AXI_READ");\n    // Packet 4645: 2 -> 11 (AXI_READ)\n    inject_packet(2, 11, 64, "AXI_READ");\n    // Packet 4646: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 4647: 7 -> 10 (AXI_WRITE)\n    inject_packet(7, 10, 64, "AXI_WRITE");\n    // Packet 4648: 12 -> 2 (AXI_WRITE)\n    inject_packet(12, 2, 64, "AXI_WRITE");\n    // Packet 4649: 13 -> 12 (AXI_WRITE)\n    inject_packet(13, 12, 64, "AXI_WRITE");\n    // Wait until cycle 958\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 958\n    // Packet 4650: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 4651: 2 -> 12 (AXI_READ)\n    inject_packet(2, 12, 64, "AXI_READ");\n    // Packet 4652: 11 -> 10 (AXI_WRITE)\n    inject_packet(11, 10, 64, "AXI_WRITE");\n    // Packet 4653: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 4654: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 959\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 959\n    // Packet 4655: 5 -> 8 (AXI_WRITE)\n    inject_packet(5, 8, 64, "AXI_WRITE");\n    // Packet 4656: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 4657: 12 -> 13 (AXI_WRITE)\n    inject_packet(12, 13, 64, "AXI_WRITE");\n    // Packet 4658: 13 -> 6 (AXI_WRITE)\n    inject_packet(13, 6, 64, "AXI_WRITE");\n    // Packet 4659: 14 -> 15 (AXI_WRITE)\n    inject_packet(14, 15, 64, "AXI_WRITE");\n    // Wait until cycle 960\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 960\n    // Packet 4660: 15 -> 3 (AXI_WRITE)\n    inject_packet(15, 3, 64, "AXI_WRITE");\n    // Wait until cycle 961\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 961\n    // Packet 4661: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 4662: 3 -> 11 (AXI_WRITE)\n    inject_packet(3, 11, 64, "AXI_WRITE");\n    // Packet 4663: 7 -> 11 (AXI_READ)\n    inject_packet(7, 11, 64, "AXI_READ");\n    // Packet 4664: 9 -> 11 (AXI_WRITE)\n    inject_packet(9, 11, 64, "AXI_WRITE");\n    // Packet 4665: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Packet 4666: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 962\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 962\n    // Packet 4667: 0 -> 8 (AXI_READ)\n    inject_packet(0, 8, 64, "AXI_READ");\n    // Packet 4668: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 4669: 9 -> 15 (AXI_READ)\n    inject_packet(9, 15, 64, "AXI_READ");\n    // Packet 4670: 11 -> 3 (AXI_READ)\n    inject_packet(11, 3, 64, "AXI_READ");\n    // Packet 4671: 13 -> 2 (AXI_WRITE)\n    inject_packet(13, 2, 64, "AXI_WRITE");\n    // Packet 4672: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Wait until cycle 963\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 963\n    // Packet 4673: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 4674: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Packet 4675: 8 -> 3 (AXI_READ)\n    inject_packet(8, 3, 64, "AXI_READ");\n    // Packet 4676: 9 -> 1 (AXI_WRITE)\n    inject_packet(9, 1, 64, "AXI_WRITE");\n    // Packet 4677: 11 -> 13 (AXI_WRITE)\n    inject_packet(11, 13, 64, "AXI_WRITE");\n    // Packet 4678: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 964\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 964\n    // Packet 4679: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 4680: 9 -> 15 (AXI_WRITE)\n    inject_packet(9, 15, 64, "AXI_WRITE");\n    // Packet 4681: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 4682: 14 -> 10 (AXI_WRITE)\n    inject_packet(14, 10, 64, "AXI_WRITE");\n    // Wait until cycle 965\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 965\n    // Packet 4683: 1 -> 8 (AXI_READ)\n    inject_packet(1, 8, 64, "AXI_READ");\n    // Packet 4684: 7 -> 5 (AXI_READ)\n    inject_packet(7, 5, 64, "AXI_READ");\n    // Packet 4685: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 4686: 10 -> 13 (AXI_READ)\n    inject_packet(10, 13, 64, "AXI_READ");\n    // Packet 4687: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Packet 4688: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Packet 4689: 15 -> 3 (AXI_READ)\n    inject_packet(15, 3, 64, "AXI_READ");\n    // Wait until cycle 966\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 966\n    // Packet 4690: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 4691: 5 -> 11 (AXI_WRITE)\n    inject_packet(5, 11, 64, "AXI_WRITE");\n    // Packet 4692: 7 -> 0 (AXI_WRITE)\n    inject_packet(7, 0, 64, "AXI_WRITE");\n    // Packet 4693: 8 -> 0 (AXI_READ)\n    inject_packet(8, 0, 64, "AXI_READ");\n    // Packet 4694: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Packet 4695: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Wait until cycle 967\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 967\n    // Packet 4696: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 4697: 7 -> 9 (AXI_WRITE)\n    inject_packet(7, 9, 64, "AXI_WRITE");\n    // Packet 4698: 12 -> 1 (AXI_READ)\n    inject_packet(12, 1, 64, "AXI_READ");\n    // Packet 4699: 13 -> 2 (AXI_READ)\n    inject_packet(13, 2, 64, "AXI_READ");\n    // Wait until cycle 968\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 968\n    // Packet 4700: 0 -> 15 (AXI_WRITE)\n    inject_packet(0, 15, 64, "AXI_WRITE");\n    // Packet 4701: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 4702: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 4703: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 4704: 12 -> 5 (AXI_WRITE)\n    inject_packet(12, 5, 64, "AXI_WRITE");\n    // Packet 4705: 13 -> 11 (AXI_READ)\n    inject_packet(13, 11, 64, "AXI_READ");\n    // Packet 4706: 15 -> 14 (AXI_READ)\n    inject_packet(15, 14, 64, "AXI_READ");\n    // Wait until cycle 969\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 969\n    // Packet 4707: 1 -> 11 (AXI_WRITE)\n    inject_packet(1, 11, 64, "AXI_WRITE");\n    // Packet 4708: 8 -> 15 (AXI_READ)\n    inject_packet(8, 15, 64, "AXI_READ");\n    // Packet 4709: 9 -> 1 (AXI_READ)\n    inject_packet(9, 1, 64, "AXI_READ");\n    // Wait until cycle 970\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 970\n    // Packet 4710: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 4711: 5 -> 7 (AXI_READ)\n    inject_packet(5, 7, 64, "AXI_READ");\n    // Packet 4712: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 4713: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 4714: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 971\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 971\n    // Packet 4715: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 4716: 1 -> 4 (AXI_READ)\n    inject_packet(1, 4, 64, "AXI_READ");\n    // Packet 4717: 3 -> 0 (AXI_WRITE)\n    inject_packet(3, 0, 64, "AXI_WRITE");\n    // Packet 4718: 9 -> 5 (AXI_WRITE)\n    inject_packet(9, 5, 64, "AXI_WRITE");\n    // Packet 4719: 10 -> 5 (AXI_READ)\n    inject_packet(10, 5, 64, "AXI_READ");\n    // Packet 4720: 14 -> 2 (AXI_WRITE)\n    inject_packet(14, 2, 64, "AXI_WRITE");\n    // Packet 4721: 15 -> 11 (AXI_READ)\n    inject_packet(15, 11, 64, "AXI_READ");\n    // Wait until cycle 972\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 972\n    // Packet 4722: 4 -> 9 (AXI_WRITE)\n    inject_packet(4, 9, 64, "AXI_WRITE");\n    // Packet 4723: 11 -> 1 (AXI_WRITE)\n    inject_packet(11, 1, 64, "AXI_WRITE");\n    // Wait until cycle 973\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 973\n    // Packet 4724: 2 -> 3 (AXI_READ)\n    inject_packet(2, 3, 64, "AXI_READ");\n    // Packet 4725: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 4726: 9 -> 6 (AXI_READ)\n    inject_packet(9, 6, 64, "AXI_READ");\n    // Packet 4727: 12 -> 14 (AXI_WRITE)\n    inject_packet(12, 14, 64, "AXI_WRITE");\n    // Packet 4728: 13 -> 3 (AXI_READ)\n    inject_packet(13, 3, 64, "AXI_READ");\n    // Wait until cycle 974\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 974\n    // Packet 4729: 3 -> 13 (AXI_WRITE)\n    inject_packet(3, 13, 64, "AXI_WRITE");\n    // Packet 4730: 5 -> 0 (AXI_READ)\n    inject_packet(5, 0, 64, "AXI_READ");\n    // Packet 4731: 10 -> 4 (AXI_READ)\n    inject_packet(10, 4, 64, "AXI_READ");\n    // Packet 4732: 13 -> 6 (AXI_READ)\n    inject_packet(13, 6, 64, "AXI_READ");\n    // Packet 4733: 14 -> 11 (AXI_READ)\n    inject_packet(14, 11, 64, "AXI_READ");\n    // Packet 4734: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 975\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 975\n    // Packet 4735: 0 -> 3 (AXI_READ)\n    inject_packet(0, 3, 64, "AXI_READ");\n    // Packet 4736: 1 -> 9 (AXI_READ)\n    inject_packet(1, 9, 64, "AXI_READ");\n    // Packet 4737: 2 -> 9 (AXI_WRITE)\n    inject_packet(2, 9, 64, "AXI_WRITE");\n    // Packet 4738: 9 -> 4 (AXI_READ)\n    inject_packet(9, 4, 64, "AXI_READ");\n    // Packet 4739: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 4740: 13 -> 15 (AXI_READ)\n    inject_packet(13, 15, 64, "AXI_READ");\n    // Wait until cycle 976\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 976\n    // Packet 4741: 1 -> 14 (AXI_WRITE)\n    inject_packet(1, 14, 64, "AXI_WRITE");\n    // Packet 4742: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 4743: 4 -> 11 (AXI_READ)\n    inject_packet(4, 11, 64, "AXI_READ");\n    // Packet 4744: 6 -> 15 (AXI_WRITE)\n    inject_packet(6, 15, 64, "AXI_WRITE");\n    // Packet 4745: 7 -> 11 (AXI_WRITE)\n    inject_packet(7, 11, 64, "AXI_WRITE");\n    // Packet 4746: 10 -> 13 (AXI_WRITE)\n    inject_packet(10, 13, 64, "AXI_WRITE");\n    // Packet 4747: 12 -> 15 (AXI_READ)\n    inject_packet(12, 15, 64, "AXI_READ");\n    // Packet 4748: 14 -> 4 (AXI_READ)\n    inject_packet(14, 4, 64, "AXI_READ");\n    // Wait until cycle 977\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 977\n    // Packet 4749: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 4750: 8 -> 7 (AXI_WRITE)\n    inject_packet(8, 7, 64, "AXI_WRITE");\n    // Packet 4751: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 4752: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Packet 4753: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Wait until cycle 978\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 978\n    // Packet 4754: 3 -> 9 (AXI_READ)\n    inject_packet(3, 9, 64, "AXI_READ");\n    // Packet 4755: 5 -> 14 (AXI_WRITE)\n    inject_packet(5, 14, 64, "AXI_WRITE");\n    // Packet 4756: 6 -> 15 (AXI_READ)\n    inject_packet(6, 15, 64, "AXI_READ");\n    // Wait until cycle 979\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 979\n    // Packet 4757: 2 -> 13 (AXI_WRITE)\n    inject_packet(2, 13, 64, "AXI_WRITE");\n    // Packet 4758: 3 -> 15 (AXI_READ)\n    inject_packet(3, 15, 64, "AXI_READ");\n    // Packet 4759: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Packet 4760: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 4761: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Wait until cycle 980\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 980\n    // Packet 4762: 1 -> 6 (AXI_READ)\n    inject_packet(1, 6, 64, "AXI_READ");\n    // Packet 4763: 3 -> 4 (AXI_WRITE)\n    inject_packet(3, 4, 64, "AXI_WRITE");\n    // Packet 4764: 5 -> 10 (AXI_READ)\n    inject_packet(5, 10, 64, "AXI_READ");\n    // Packet 4765: 6 -> 3 (AXI_READ)\n    inject_packet(6, 3, 64, "AXI_READ");\n    // Packet 4766: 8 -> 12 (AXI_WRITE)\n    inject_packet(8, 12, 64, "AXI_WRITE");\n    // Packet 4767: 10 -> 9 (AXI_WRITE)\n    inject_packet(10, 9, 64, "AXI_WRITE");\n    // Packet 4768: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Wait until cycle 981\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 981\n    // Packet 4769: 1 -> 5 (AXI_READ)\n    inject_packet(1, 5, 64, "AXI_READ");\n    // Packet 4770: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 4771: 3 -> 5 (AXI_READ)\n    inject_packet(3, 5, 64, "AXI_READ");\n    // Packet 4772: 5 -> 8 (AXI_READ)\n    inject_packet(5, 8, 64, "AXI_READ");\n    // Packet 4773: 11 -> 8 (AXI_WRITE)\n    inject_packet(11, 8, 64, "AXI_WRITE");\n    // Packet 4774: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 982\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 982\n    // Packet 4775: 2 -> 3 (AXI_WRITE)\n    inject_packet(2, 3, 64, "AXI_WRITE");\n    // Packet 4776: 4 -> 13 (AXI_READ)\n    inject_packet(4, 13, 64, "AXI_READ");\n    // Packet 4777: 5 -> 2 (AXI_WRITE)\n    inject_packet(5, 2, 64, "AXI_WRITE");\n    // Packet 4778: 7 -> 2 (AXI_READ)\n    inject_packet(7, 2, 64, "AXI_READ");\n    // Packet 4779: 13 -> 4 (AXI_READ)\n    inject_packet(13, 4, 64, "AXI_READ");\n    // Packet 4780: 15 -> 6 (AXI_WRITE)\n    inject_packet(15, 6, 64, "AXI_WRITE");\n    // Wait until cycle 983\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 983\n    // Packet 4781: 0 -> 15 (AXI_READ)\n    inject_packet(0, 15, 64, "AXI_READ");\n    // Packet 4782: 2 -> 5 (AXI_READ)\n    inject_packet(2, 5, 64, "AXI_READ");\n    // Packet 4783: 5 -> 1 (AXI_WRITE)\n    inject_packet(5, 1, 64, "AXI_WRITE");\n    // Packet 4784: 8 -> 1 (AXI_WRITE)\n    inject_packet(8, 1, 64, "AXI_WRITE");\n    // Packet 4785: 13 -> 14 (AXI_READ)\n    inject_packet(13, 14, 64, "AXI_READ");\n    // Wait until cycle 984\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 984\n    // Packet 4786: 3 -> 4 (AXI_READ)\n    inject_packet(3, 4, 64, "AXI_READ");\n    // Packet 4787: 8 -> 2 (AXI_READ)\n    inject_packet(8, 2, 64, "AXI_READ");\n    // Packet 4788: 11 -> 9 (AXI_READ)\n    inject_packet(11, 9, 64, "AXI_READ");\n    // Packet 4789: 13 -> 9 (AXI_READ)\n    inject_packet(13, 9, 64, "AXI_READ");\n    // Wait until cycle 985\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 985\n    // Packet 4790: 1 -> 11 (AXI_READ)\n    inject_packet(1, 11, 64, "AXI_READ");\n    // Packet 4791: 2 -> 10 (AXI_WRITE)\n    inject_packet(2, 10, 64, "AXI_WRITE");\n    // Packet 4792: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 4793: 9 -> 12 (AXI_WRITE)\n    inject_packet(9, 12, 64, "AXI_WRITE");\n    // Packet 4794: 12 -> 7 (AXI_READ)\n    inject_packet(12, 7, 64, "AXI_READ");\n    // Packet 4795: 13 -> 4 (AXI_WRITE)\n    inject_packet(13, 4, 64, "AXI_WRITE");\n    // Wait until cycle 986\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 986\n    // Packet 4796: 0 -> 4 (AXI_READ)\n    inject_packet(0, 4, 64, "AXI_READ");\n    // Packet 4797: 6 -> 5 (AXI_WRITE)\n    inject_packet(6, 5, 64, "AXI_WRITE");\n    // Packet 4798: 7 -> 12 (AXI_WRITE)\n    inject_packet(7, 12, 64, "AXI_WRITE");\n    // Packet 4799: 11 -> 4 (AXI_WRITE)\n    inject_packet(11, 4, 64, "AXI_WRITE");\n    // Packet 4800: 12 -> 9 (AXI_READ)\n    inject_packet(12, 9, 64, "AXI_READ");\n    // Wait until cycle 987\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 987\n    // Packet 4801: 3 -> 2 (AXI_WRITE)\n    inject_packet(3, 2, 64, "AXI_WRITE");\n    // Packet 4802: 6 -> 0 (AXI_READ)\n    inject_packet(6, 0, 64, "AXI_READ");\n    // Packet 4803: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 4804: 14 -> 3 (AXI_READ)\n    inject_packet(14, 3, 64, "AXI_READ");\n    // Wait until cycle 988\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 988\n    // Packet 4805: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 4806: 8 -> 11 (AXI_WRITE)\n    inject_packet(8, 11, 64, "AXI_WRITE");\n    // Packet 4807: 9 -> 5 (AXI_READ)\n    inject_packet(9, 5, 64, "AXI_READ");\n    // Packet 4808: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 4809: 13 -> 8 (AXI_WRITE)\n    inject_packet(13, 8, 64, "AXI_WRITE");\n    // Wait until cycle 989\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 989\n    // Packet 4810: 0 -> 5 (AXI_READ)\n    inject_packet(0, 5, 64, "AXI_READ");\n    // Packet 4811: 2 -> 0 (AXI_READ)\n    inject_packet(2, 0, 64, "AXI_READ");\n    // Packet 4812: 4 -> 14 (AXI_WRITE)\n    inject_packet(4, 14, 64, "AXI_WRITE");\n    // Packet 4813: 6 -> 13 (AXI_READ)\n    inject_packet(6, 13, 64, "AXI_READ");\n    // Packet 4814: 9 -> 2 (AXI_WRITE)\n    inject_packet(9, 2, 64, "AXI_WRITE");\n    // Packet 4815: 15 -> 7 (AXI_WRITE)\n    inject_packet(15, 7, 64, "AXI_WRITE");\n    // Wait until cycle 990\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 990\n    // Packet 4816: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 4817: 4 -> 6 (AXI_READ)\n    inject_packet(4, 6, 64, "AXI_READ");\n    // Packet 4818: 6 -> 1 (AXI_READ)\n    inject_packet(6, 1, 64, "AXI_READ");\n    // Packet 4819: 9 -> 6 (AXI_WRITE)\n    inject_packet(9, 6, 64, "AXI_WRITE");\n    // Packet 4820: 10 -> 6 (AXI_WRITE)\n    inject_packet(10, 6, 64, "AXI_WRITE");\n    // Packet 4821: 11 -> 6 (AXI_WRITE)\n    inject_packet(11, 6, 64, "AXI_WRITE");\n    // Wait until cycle 991\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 991\n    // Packet 4822: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Wait until cycle 992\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 992\n    // Packet 4823: 0 -> 5 (AXI_WRITE)\n    inject_packet(0, 5, 64, "AXI_WRITE");\n    // Packet 4824: 3 -> 7 (AXI_READ)\n    inject_packet(3, 7, 64, "AXI_READ");\n    // Packet 4825: 12 -> 10 (AXI_READ)\n    inject_packet(12, 10, 64, "AXI_READ");\n    // Wait until cycle 993\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 993\n    // Packet 4826: 2 -> 4 (AXI_WRITE)\n    inject_packet(2, 4, 64, "AXI_WRITE");\n    // Packet 4827: 6 -> 11 (AXI_WRITE)\n    inject_packet(6, 11, 64, "AXI_WRITE");\n    // Packet 4828: 8 -> 10 (AXI_READ)\n    inject_packet(8, 10, 64, "AXI_READ");\n    // Packet 4829: 13 -> 12 (AXI_READ)\n    inject_packet(13, 12, 64, "AXI_READ");\n    // Packet 4830: 14 -> 7 (AXI_WRITE)\n    inject_packet(14, 7, 64, "AXI_WRITE");\n    // Wait until cycle 994\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 994\n    // Packet 4831: 4 -> 15 (AXI_WRITE)\n    inject_packet(4, 15, 64, "AXI_WRITE");\n    // Packet 4832: 11 -> 10 (AXI_READ)\n    inject_packet(11, 10, 64, "AXI_READ");\n    // Packet 4833: 13 -> 10 (AXI_READ)\n    inject_packet(13, 10, 64, "AXI_READ");\n    // Packet 4834: 14 -> 7 (AXI_READ)\n    inject_packet(14, 7, 64, "AXI_READ");\n    // Wait until cycle 995\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 995\n    // Packet 4835: 0 -> 11 (AXI_READ)\n    inject_packet(0, 11, 64, "AXI_READ");\n    // Packet 4836: 4 -> 1 (AXI_WRITE)\n    inject_packet(4, 1, 64, "AXI_WRITE");\n    // Packet 4837: 10 -> 2 (AXI_WRITE)\n    inject_packet(10, 2, 64, "AXI_WRITE");\n    // Packet 4838: 11 -> 1 (AXI_READ)\n    inject_packet(11, 1, 64, "AXI_READ");\n    // Packet 4839: 15 -> 13 (AXI_READ)\n    inject_packet(15, 13, 64, "AXI_READ");\n    // Wait until cycle 996\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 996\n    // Packet 4840: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 4841: 7 -> 13 (AXI_READ)\n    inject_packet(7, 13, 64, "AXI_READ");\n    // Packet 4842: 11 -> 13 (AXI_READ)\n    inject_packet(11, 13, 64, "AXI_READ");\n    // Wait until cycle 997\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 997\n    // Packet 4843: 1 -> 4 (AXI_WRITE)\n    inject_packet(1, 4, 64, "AXI_WRITE");\n    // Packet 4844: 2 -> 6 (AXI_WRITE)\n    inject_packet(2, 6, 64, "AXI_WRITE");\n    // Packet 4845: 4 -> 7 (AXI_READ)\n    inject_packet(4, 7, 64, "AXI_READ");\n    // Packet 4846: 5 -> 6 (AXI_WRITE)\n    inject_packet(5, 6, 64, "AXI_WRITE");\n    // Packet 4847: 6 -> 12 (AXI_READ)\n    inject_packet(6, 12, 64, "AXI_READ");\n    // Packet 4848: 7 -> 3 (AXI_READ)\n    inject_packet(7, 3, 64, "AXI_READ");\n    // Packet 4849: 8 -> 5 (AXI_READ)\n    inject_packet(8, 5, 64, "AXI_READ");\n    // Packet 4850: 15 -> 14 (AXI_WRITE)\n    inject_packet(15, 14, 64, "AXI_WRITE");\n    // Wait until cycle 998\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 998\n    // Packet 4851: 0 -> 2 (AXI_WRITE)\n    inject_packet(0, 2, 64, "AXI_WRITE");\n    // Packet 4852: 7 -> 9 (AXI_READ)\n    inject_packet(7, 9, 64, "AXI_READ");\n    // Packet 4853: 8 -> 11 (AXI_READ)\n    inject_packet(8, 11, 64, "AXI_READ");\n    // Packet 4854: 9 -> 0 (AXI_WRITE)\n    inject_packet(9, 0, 64, "AXI_WRITE");\n    // Packet 4855: 10 -> 5 (AXI_WRITE)\n    inject_packet(10, 5, 64, "AXI_WRITE");\n    // Packet 4856: 13 -> 3 (AXI_WRITE)\n    inject_packet(13, 3, 64, "AXI_WRITE");\n    // Packet 4857: 14 -> 10 (AXI_READ)\n    inject_packet(14, 10, 64, "AXI_READ");\n    // Packet 4858: 15 -> 10 (AXI_READ)\n    inject_packet(15, 10, 64, "AXI_READ");\n    // Wait until cycle 999\n    repeat(1) @(posedge clk);\n    // Inject packets at cycle 999\n    // Packet 4859: 3 -> 0 (AXI_READ)\n    inject_packet(3, 0, 64, "AXI_READ");\n    // Packet 4860: 4 -> 7 (AXI_WRITE)\n    inject_packet(4, 7, 64, "AXI_WRITE");\n    // Packet 4861: 10 -> 15 (AXI_READ)\n    inject_packet(10, 15, 64, "AXI_READ");\n    // Packet 4862: 11 -> 7 (AXI_READ)\n    inject_packet(11, 7, 64, "AXI_READ");\n
    // Wait for completion
    repeat(1000) @(posedge clk);
    
    $display("Traffic pattern simulation completed");
    $finish;
  end
  
  task inject_packet(
    input int src_node,
    input int dst_node, 
    input int size_bytes,
    input string pkt_type
  );
    // Implementation depends on specific interface
    $display("[%0t] Injecting %s packet: %0d -> %0d (%0d bytes)", 
             $time, pkt_type, src_node, dst_node, size_bytes);
  endtask

endmodule
