`timescale 1ns / 1ps

module tb_nebula_top_traffic;
    import nebula_pkg::*;

    // Parameters
    parameter int MESH_WIDTH = 4;
    parameter int MESH_HEIGHT = 4;
    parameter int NUM_NODES = 16;
    parameter int CONFIG_ADDR_WIDTH = 16;
    parameter int CONFIG_DATA_WIDTH = 32;
    parameter bit ENABLE_AXI = 1'b1;
    parameter bit ENABLE_CHI = 1'b1;
    parameter bit ENABLE_PERFORMANCE_MONITORING = 1'b1;

    // Traffic data type definition
    typedef struct {
        int timestamp;
        int source_node;
        int dest_node;
        string packet_type;
        int size_bytes;
    } traffic_entry_t;
    
    parameter int TRAFFIC_SIZE = 1581;
    traffic_entry_t traffic_data[TRAFFIC_SIZE];

    // Clock and reset
    logic clk;
    logic rst_n;
    
    // System Configuration Interface  
    logic                           config_req_valid;
    logic                           config_req_ready;
    logic [CONFIG_ADDR_WIDTH-1:0]  config_req_addr;
    logic [CONFIG_DATA_WIDTH-1:0]  config_req_data;
    logic                           config_req_write;
    logic                           config_resp_valid;
    logic                           config_resp_ready;
    logic [CONFIG_DATA_WIDTH-1:0]  config_resp_data;
    logic                           config_resp_error;
    
    // Memory interfaces
    logic [NUM_NODES-1:0]                     mem_req_valid;
    logic [NUM_NODES-1:0]                     mem_req_ready;
    logic [NUM_NODES-1:0][CHI_REQ_ADDR_WIDTH-1:0] mem_req_addr;
    logic [NUM_NODES-1:0]                     mem_req_write;
    logic [NUM_NODES-1:0][CHI_DATA_WIDTH-1:0] mem_req_data;
    logic [NUM_NODES-1:0][CHI_BE_WIDTH-1:0]   mem_req_be;
    logic [NUM_NODES-1:0]                     mem_resp_valid;
    logic [NUM_NODES-1:0]                     mem_resp_ready;
    logic [NUM_NODES-1:0][CHI_DATA_WIDTH-1:0] mem_resp_data;
    logic [NUM_NODES-1:0]                     mem_resp_error;
    
    // AXI interfaces  
    logic [NUM_NODES-1:0]                     axi_aw_valid;
    logic [NUM_NODES-1:0]                     axi_aw_ready;
    axi_aw_t [NUM_NODES-1:0]                  axi_aw;
    logic [NUM_NODES-1:0]                     axi_w_valid;
    logic [NUM_NODES-1:0]                     axi_w_ready;
    axi_w_t [NUM_NODES-1:0]                   axi_w;
    logic [NUM_NODES-1:0]                     axi_b_valid;
    logic [NUM_NODES-1:0]                     axi_b_ready;
    axi_b_t [NUM_NODES-1:0]                   axi_b;
    logic [NUM_NODES-1:0]                     axi_ar_valid;
    logic [NUM_NODES-1:0]                     axi_ar_ready;
    axi_ar_t [NUM_NODES-1:0]                  axi_ar;
    logic [NUM_NODES-1:0]                     axi_r_valid;
    logic [NUM_NODES-1:0]                     axi_r_ready;
    axi_r_t [NUM_NODES-1:0]                   axi_r;
    
    // CHI interfaces
    logic [NUM_NODES-1:0]                     chi_req_valid;
    logic [NUM_NODES-1:0]                     chi_req_ready;
    chi_req_t [NUM_NODES-1:0]                 chi_req;
    logic [NUM_NODES-1:0]                     chi_resp_valid;
    logic [NUM_NODES-1:0]                     chi_resp_ready;
    chi_resp_t [NUM_NODES-1:0]                chi_resp;
    logic [NUM_NODES-1:0]                     chi_dat_req_valid;
    logic [NUM_NODES-1:0]                     chi_dat_req_ready;
    chi_data_t [NUM_NODES-1:0]                chi_dat_req;
    logic [NUM_NODES-1:0]                     chi_dat_resp_valid;
    logic [NUM_NODES-1:0]                     chi_dat_resp_ready;
    chi_data_t [NUM_NODES-1:0]                chi_dat_resp;
    
    // System Status and Debug  
    logic [31:0]                              system_status;
    logic [31:0]                              error_status;
    logic [31:0]                              performance_counters [15:0];
    logic                                     debug_trace_valid;
    logic [63:0]                             debug_trace_data;
    logic [7:0]                              debug_trace_node_id;

    // DUT instantiation
    nebula_top #(
        .MESH_WIDTH(MESH_WIDTH),
        .MESH_HEIGHT(MESH_HEIGHT),
        .NUM_NODES(NUM_NODES),
        .CONFIG_ADDR_WIDTH(CONFIG_ADDR_WIDTH),
        .CONFIG_DATA_WIDTH(CONFIG_DATA_WIDTH),
        .ENABLE_AXI(ENABLE_AXI),
        .ENABLE_CHI(ENABLE_CHI),
        .ENABLE_PERFORMANCE_MONITORING(ENABLE_PERFORMANCE_MONITORING)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .config_req_valid(config_req_valid),
        .config_req_ready(config_req_ready),
        .config_req_addr(config_req_addr),
        .config_req_data(config_req_data),
        .config_req_write(config_req_write),
        .config_resp_valid(config_resp_valid),
        .config_resp_ready(config_resp_ready),
        .config_resp_data(config_resp_data),
        .config_resp_error(config_resp_error),
        .mem_req_valid(mem_req_valid),
        .mem_req_ready(mem_req_ready),
        .mem_req_addr(mem_req_addr),   
        .mem_req_write(mem_req_write),
        .mem_req_data(mem_req_data),
        .mem_req_be(mem_req_be),
        .mem_resp_valid(mem_resp_valid),   
        .mem_resp_ready(mem_resp_ready),
        .mem_resp_data(mem_resp_data),
        .mem_resp_error(mem_resp_error),
        .axi_aw_valid(axi_aw_valid),   
        .axi_aw_ready(axi_aw_ready),
        .axi_aw(axi_aw),
        .axi_w_valid(axi_w_valid),    
        .axi_w_ready(axi_w_ready),
        .axi_w(axi_w),    
        .axi_b_valid(axi_b_valid),    
        .axi_b_ready(axi_b_ready),
        .axi_b(axi_b),    
        .axi_ar_valid(axi_ar_valid),   
        .axi_ar_ready(axi_ar_ready),
        .axi_ar(axi_ar),   
        .axi_r_valid(axi_r_valid),    
        .axi_r_ready(axi_r_ready),
        .axi_r(axi_r),    
        .chi_req_valid(chi_req_valid),     
        .chi_req_ready(chi_req_ready),
        .chi_req(chi_req),
        .chi_resp_valid(chi_resp_valid),
        .chi_resp_ready(chi_resp_ready),
        .chi_resp(chi_resp),
        .chi_dat_req_valid(chi_dat_req_valid),
        .chi_dat_req_ready(chi_dat_req_ready),
        .chi_dat_req(chi_dat_req),
        .chi_dat_resp_valid(chi_dat_resp_valid),
        .chi_dat_resp_ready(chi_dat_resp_ready),
        .chi_dat_resp(chi_dat_resp),
        .system_status(system_status),
        .error_status(error_status),
        .performance_counters(performance_counters),
        .debug_trace_valid(debug_trace_valid),
        .debug_trace_node_id(debug_trace_node_id),
        .debug_trace_data(debug_trace_data)
    );
    
    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 100MHz clock
    end
    
    // Reset and test sequence
    initial begin
        // Initialize signals
        rst_n = 0;
        config_req_valid = 0;
        config_req_addr = 0;
        config_req_data = 0;
        config_req_write = 0;
        config_resp_ready = 1;
        
        // Initialize memory interfaces
        mem_req_ready = '1;
        mem_resp_valid = '0;
        mem_resp_data = '0;
        mem_resp_error = '0;
        
        // Initialize AXI interfaces
        axi_aw_valid = '0;
        axi_aw = '0;
        axi_w_valid = '0;
        axi_w = '0;
        axi_b_ready = '1;
        axi_ar_valid = '0;
        axi_ar = '0;
        axi_r_ready = '1;
        
        // Initialize CHI interfaces
        chi_req_valid = '0;
        chi_req = '0;
        chi_resp_ready = '1;
        chi_dat_req_valid = '0;
        chi_dat_req = '0;
        chi_dat_resp_ready = '1;
        
        // Apply reset
        #20;
        rst_n = 1;
        #20;
        
        $display("🔧 Starting NoC traffic simulation with %0d nodes...", NUM_NODES);
        $display("🔧 Traffic size: %0d entries", TRAFFIC_SIZE);
        
        // Wait for system to stabilize
        repeat(100) @(posedge clk);
        $display("🔧 System stabilization complete");
        
        // Enable VCD dumping
        $dumpfile("tb_nebula_traffic.vcd");
        $dumpvars(0, tb_nebula_top_traffic);
        $display("🔧 VCD dumping enabled");
        
        // Load traffic data
        $display("📝 Loading traffic data...");
        traffic_data[0].timestamp = 0;
        traffic_data[0].source_node = 1;
        traffic_data[0].dest_node = 5;
        traffic_data[0].packet_type = "AXI_WRITE";
        traffic_data[0].size_bytes = 64;
        traffic_data[1].timestamp = 0;
        traffic_data[1].source_node = 6;
        traffic_data[1].dest_node = 7;
        traffic_data[1].packet_type = "AXI_READ";
        traffic_data[1].size_bytes = 64;
        traffic_data[2].timestamp = 0;
        traffic_data[2].source_node = 7;
        traffic_data[2].dest_node = 3;
        traffic_data[2].packet_type = "AXI_WRITE";
        traffic_data[2].size_bytes = 64;
        traffic_data[3].timestamp = 0;
        traffic_data[3].source_node = 9;
        traffic_data[3].dest_node = 3;
        traffic_data[3].packet_type = "CHI_WRITE";
        traffic_data[3].size_bytes = 64;
        traffic_data[4].timestamp = 0;
        traffic_data[4].source_node = 13;
        traffic_data[4].dest_node = 12;
        traffic_data[4].packet_type = "AXI_WRITE";
        traffic_data[4].size_bytes = 64;
        traffic_data[5].timestamp = 1;
        traffic_data[5].source_node = 3;
        traffic_data[5].dest_node = 1;
        traffic_data[5].packet_type = "CHI_READ";
        traffic_data[5].size_bytes = 64;
        traffic_data[6].timestamp = 2;
        traffic_data[6].source_node = 1;
        traffic_data[6].dest_node = 4;
        traffic_data[6].packet_type = "CHI_READ";
        traffic_data[6].size_bytes = 64;
        traffic_data[7].timestamp = 2;
        traffic_data[7].source_node = 13;
        traffic_data[7].dest_node = 10;
        traffic_data[7].packet_type = "AXI_WRITE";
        traffic_data[7].size_bytes = 64;
        traffic_data[8].timestamp = 3;
        traffic_data[8].source_node = 7;
        traffic_data[8].dest_node = 14;
        traffic_data[8].packet_type = "AXI_READ";
        traffic_data[8].size_bytes = 64;
        traffic_data[9].timestamp = 3;
        traffic_data[9].source_node = 10;
        traffic_data[9].dest_node = 15;
        traffic_data[9].packet_type = "CHI_READ";
        traffic_data[9].size_bytes = 64;
        traffic_data[10].timestamp = 5;
        traffic_data[10].source_node = 14;
        traffic_data[10].dest_node = 11;
        traffic_data[10].packet_type = "CHI_READ";
        traffic_data[10].size_bytes = 64;
        traffic_data[11].timestamp = 7;
        traffic_data[11].source_node = 5;
        traffic_data[11].dest_node = 12;
        traffic_data[11].packet_type = "CHI_WRITE";
        traffic_data[11].size_bytes = 64;
        traffic_data[12].timestamp = 8;
        traffic_data[12].source_node = 10;
        traffic_data[12].dest_node = 0;
        traffic_data[12].packet_type = "AXI_WRITE";
        traffic_data[12].size_bytes = 64;
        traffic_data[13].timestamp = 8;
        traffic_data[13].source_node = 12;
        traffic_data[13].dest_node = 11;
        traffic_data[13].packet_type = "AXI_READ";
        traffic_data[13].size_bytes = 64;
        traffic_data[14].timestamp = 9;
        traffic_data[14].source_node = 0;
        traffic_data[14].dest_node = 4;
        traffic_data[14].packet_type = "CHI_READ";
        traffic_data[14].size_bytes = 64;
        traffic_data[15].timestamp = 9;
        traffic_data[15].source_node = 10;
        traffic_data[15].dest_node = 6;
        traffic_data[15].packet_type = "CHI_READ";
        traffic_data[15].size_bytes = 64;
        traffic_data[16].timestamp = 10;
        traffic_data[16].source_node = 0;
        traffic_data[16].dest_node = 7;
        traffic_data[16].packet_type = "CHI_READ";
        traffic_data[16].size_bytes = 64;
        traffic_data[17].timestamp = 10;
        traffic_data[17].source_node = 9;
        traffic_data[17].dest_node = 13;
        traffic_data[17].packet_type = "AXI_READ";
        traffic_data[17].size_bytes = 64;
        traffic_data[18].timestamp = 10;
        traffic_data[18].source_node = 10;
        traffic_data[18].dest_node = 8;
        traffic_data[18].packet_type = "AXI_READ";
        traffic_data[18].size_bytes = 64;
        traffic_data[19].timestamp = 11;
        traffic_data[19].source_node = 2;
        traffic_data[19].dest_node = 7;
        traffic_data[19].packet_type = "AXI_READ";
        traffic_data[19].size_bytes = 64;
        traffic_data[20].timestamp = 12;
        traffic_data[20].source_node = 2;
        traffic_data[20].dest_node = 10;
        traffic_data[20].packet_type = "CHI_WRITE";
        traffic_data[20].size_bytes = 64;
        traffic_data[21].timestamp = 12;
        traffic_data[21].source_node = 7;
        traffic_data[21].dest_node = 2;
        traffic_data[21].packet_type = "AXI_READ";
        traffic_data[21].size_bytes = 64;
        traffic_data[22].timestamp = 13;
        traffic_data[22].source_node = 12;
        traffic_data[22].dest_node = 7;
        traffic_data[22].packet_type = "AXI_READ";
        traffic_data[22].size_bytes = 64;
        traffic_data[23].timestamp = 13;
        traffic_data[23].source_node = 13;
        traffic_data[23].dest_node = 3;
        traffic_data[23].packet_type = "CHI_READ";
        traffic_data[23].size_bytes = 64;
        traffic_data[24].timestamp = 14;
        traffic_data[24].source_node = 0;
        traffic_data[24].dest_node = 4;
        traffic_data[24].packet_type = "CHI_READ";
        traffic_data[24].size_bytes = 64;
        traffic_data[25].timestamp = 15;
        traffic_data[25].source_node = 9;
        traffic_data[25].dest_node = 11;
        traffic_data[25].packet_type = "CHI_WRITE";
        traffic_data[25].size_bytes = 64;
        traffic_data[26].timestamp = 15;
        traffic_data[26].source_node = 11;
        traffic_data[26].dest_node = 5;
        traffic_data[26].packet_type = "AXI_WRITE";
        traffic_data[26].size_bytes = 64;
        traffic_data[27].timestamp = 16;
        traffic_data[27].source_node = 1;
        traffic_data[27].dest_node = 2;
        traffic_data[27].packet_type = "AXI_WRITE";
        traffic_data[27].size_bytes = 64;
        traffic_data[28].timestamp = 17;
        traffic_data[28].source_node = 9;
        traffic_data[28].dest_node = 12;
        traffic_data[28].packet_type = "CHI_READ";
        traffic_data[28].size_bytes = 64;
        traffic_data[29].timestamp = 18;
        traffic_data[29].source_node = 2;
        traffic_data[29].dest_node = 8;
        traffic_data[29].packet_type = "AXI_WRITE";
        traffic_data[29].size_bytes = 64;
        traffic_data[30].timestamp = 18;
        traffic_data[30].source_node = 12;
        traffic_data[30].dest_node = 13;
        traffic_data[30].packet_type = "CHI_READ";
        traffic_data[30].size_bytes = 64;
        traffic_data[31].timestamp = 19;
        traffic_data[31].source_node = 2;
        traffic_data[31].dest_node = 15;
        traffic_data[31].packet_type = "CHI_READ";
        traffic_data[31].size_bytes = 64;
        traffic_data[32].timestamp = 20;
        traffic_data[32].source_node = 0;
        traffic_data[32].dest_node = 15;
        traffic_data[32].packet_type = "AXI_WRITE";
        traffic_data[32].size_bytes = 64;
        traffic_data[33].timestamp = 20;
        traffic_data[33].source_node = 2;
        traffic_data[33].dest_node = 11;
        traffic_data[33].packet_type = "CHI_READ";
        traffic_data[33].size_bytes = 64;
        traffic_data[34].timestamp = 22;
        traffic_data[34].source_node = 3;
        traffic_data[34].dest_node = 13;
        traffic_data[34].packet_type = "AXI_WRITE";
        traffic_data[34].size_bytes = 64;
        traffic_data[35].timestamp = 22;
        traffic_data[35].source_node = 7;
        traffic_data[35].dest_node = 3;
        traffic_data[35].packet_type = "CHI_WRITE";
        traffic_data[35].size_bytes = 64;
        traffic_data[36].timestamp = 25;
        traffic_data[36].source_node = 7;
        traffic_data[36].dest_node = 2;
        traffic_data[36].packet_type = "AXI_WRITE";
        traffic_data[36].size_bytes = 64;
        traffic_data[37].timestamp = 25;
        traffic_data[37].source_node = 14;
        traffic_data[37].dest_node = 13;
        traffic_data[37].packet_type = "CHI_WRITE";
        traffic_data[37].size_bytes = 64;
        traffic_data[38].timestamp = 26;
        traffic_data[38].source_node = 2;
        traffic_data[38].dest_node = 15;
        traffic_data[38].packet_type = "CHI_WRITE";
        traffic_data[38].size_bytes = 64;
        traffic_data[39].timestamp = 27;
        traffic_data[39].source_node = 11;
        traffic_data[39].dest_node = 6;
        traffic_data[39].packet_type = "AXI_WRITE";
        traffic_data[39].size_bytes = 64;
        traffic_data[40].timestamp = 28;
        traffic_data[40].source_node = 9;
        traffic_data[40].dest_node = 5;
        traffic_data[40].packet_type = "AXI_WRITE";
        traffic_data[40].size_bytes = 64;
        traffic_data[41].timestamp = 29;
        traffic_data[41].source_node = 0;
        traffic_data[41].dest_node = 3;
        traffic_data[41].packet_type = "AXI_WRITE";
        traffic_data[41].size_bytes = 64;
        traffic_data[42].timestamp = 29;
        traffic_data[42].source_node = 14;
        traffic_data[42].dest_node = 4;
        traffic_data[42].packet_type = "CHI_WRITE";
        traffic_data[42].size_bytes = 64;
        traffic_data[43].timestamp = 30;
        traffic_data[43].source_node = 1;
        traffic_data[43].dest_node = 12;
        traffic_data[43].packet_type = "AXI_WRITE";
        traffic_data[43].size_bytes = 64;
        traffic_data[44].timestamp = 32;
        traffic_data[44].source_node = 1;
        traffic_data[44].dest_node = 15;
        traffic_data[44].packet_type = "CHI_WRITE";
        traffic_data[44].size_bytes = 64;
        traffic_data[45].timestamp = 32;
        traffic_data[45].source_node = 6;
        traffic_data[45].dest_node = 14;
        traffic_data[45].packet_type = "CHI_READ";
        traffic_data[45].size_bytes = 64;
        traffic_data[46].timestamp = 32;
        traffic_data[46].source_node = 14;
        traffic_data[46].dest_node = 3;
        traffic_data[46].packet_type = "AXI_READ";
        traffic_data[46].size_bytes = 64;
        traffic_data[47].timestamp = 33;
        traffic_data[47].source_node = 6;
        traffic_data[47].dest_node = 4;
        traffic_data[47].packet_type = "AXI_WRITE";
        traffic_data[47].size_bytes = 64;
        traffic_data[48].timestamp = 35;
        traffic_data[48].source_node = 5;
        traffic_data[48].dest_node = 0;
        traffic_data[48].packet_type = "CHI_READ";
        traffic_data[48].size_bytes = 64;
        traffic_data[49].timestamp = 35;
        traffic_data[49].source_node = 15;
        traffic_data[49].dest_node = 13;
        traffic_data[49].packet_type = "CHI_WRITE";
        traffic_data[49].size_bytes = 64;
        traffic_data[50].timestamp = 36;
        traffic_data[50].source_node = 1;
        traffic_data[50].dest_node = 8;
        traffic_data[50].packet_type = "AXI_READ";
        traffic_data[50].size_bytes = 64;
        traffic_data[51].timestamp = 36;
        traffic_data[51].source_node = 7;
        traffic_data[51].dest_node = 3;
        traffic_data[51].packet_type = "AXI_READ";
        traffic_data[51].size_bytes = 64;
        traffic_data[52].timestamp = 37;
        traffic_data[52].source_node = 3;
        traffic_data[52].dest_node = 12;
        traffic_data[52].packet_type = "AXI_READ";
        traffic_data[52].size_bytes = 64;
        traffic_data[53].timestamp = 37;
        traffic_data[53].source_node = 10;
        traffic_data[53].dest_node = 0;
        traffic_data[53].packet_type = "CHI_WRITE";
        traffic_data[53].size_bytes = 64;
        traffic_data[54].timestamp = 38;
        traffic_data[54].source_node = 13;
        traffic_data[54].dest_node = 2;
        traffic_data[54].packet_type = "CHI_READ";
        traffic_data[54].size_bytes = 64;
        traffic_data[55].timestamp = 39;
        traffic_data[55].source_node = 12;
        traffic_data[55].dest_node = 3;
        traffic_data[55].packet_type = "AXI_READ";
        traffic_data[55].size_bytes = 64;
        traffic_data[56].timestamp = 40;
        traffic_data[56].source_node = 0;
        traffic_data[56].dest_node = 13;
        traffic_data[56].packet_type = "AXI_WRITE";
        traffic_data[56].size_bytes = 64;
        traffic_data[57].timestamp = 40;
        traffic_data[57].source_node = 8;
        traffic_data[57].dest_node = 5;
        traffic_data[57].packet_type = "CHI_WRITE";
        traffic_data[57].size_bytes = 64;
        traffic_data[58].timestamp = 42;
        traffic_data[58].source_node = 13;
        traffic_data[58].dest_node = 14;
        traffic_data[58].packet_type = "AXI_READ";
        traffic_data[58].size_bytes = 64;
        traffic_data[59].timestamp = 45;
        traffic_data[59].source_node = 5;
        traffic_data[59].dest_node = 12;
        traffic_data[59].packet_type = "CHI_WRITE";
        traffic_data[59].size_bytes = 64;
        traffic_data[60].timestamp = 45;
        traffic_data[60].source_node = 13;
        traffic_data[60].dest_node = 8;
        traffic_data[60].packet_type = "CHI_READ";
        traffic_data[60].size_bytes = 64;
        traffic_data[61].timestamp = 47;
        traffic_data[61].source_node = 4;
        traffic_data[61].dest_node = 1;
        traffic_data[61].packet_type = "AXI_WRITE";
        traffic_data[61].size_bytes = 64;
        traffic_data[62].timestamp = 47;
        traffic_data[62].source_node = 10;
        traffic_data[62].dest_node = 11;
        traffic_data[62].packet_type = "AXI_READ";
        traffic_data[62].size_bytes = 64;
        traffic_data[63].timestamp = 47;
        traffic_data[63].source_node = 14;
        traffic_data[63].dest_node = 12;
        traffic_data[63].packet_type = "AXI_READ";
        traffic_data[63].size_bytes = 64;
        traffic_data[64].timestamp = 48;
        traffic_data[64].source_node = 6;
        traffic_data[64].dest_node = 14;
        traffic_data[64].packet_type = "CHI_WRITE";
        traffic_data[64].size_bytes = 64;
        traffic_data[65].timestamp = 48;
        traffic_data[65].source_node = 14;
        traffic_data[65].dest_node = 12;
        traffic_data[65].packet_type = "CHI_WRITE";
        traffic_data[65].size_bytes = 64;
        traffic_data[66].timestamp = 50;
        traffic_data[66].source_node = 7;
        traffic_data[66].dest_node = 10;
        traffic_data[66].packet_type = "CHI_WRITE";
        traffic_data[66].size_bytes = 64;
        traffic_data[67].timestamp = 51;
        traffic_data[67].source_node = 4;
        traffic_data[67].dest_node = 11;
        traffic_data[67].packet_type = "AXI_READ";
        traffic_data[67].size_bytes = 64;
        traffic_data[68].timestamp = 51;
        traffic_data[68].source_node = 9;
        traffic_data[68].dest_node = 4;
        traffic_data[68].packet_type = "CHI_READ";
        traffic_data[68].size_bytes = 64;
        traffic_data[69].timestamp = 53;
        traffic_data[69].source_node = 3;
        traffic_data[69].dest_node = 9;
        traffic_data[69].packet_type = "AXI_READ";
        traffic_data[69].size_bytes = 64;
        traffic_data[70].timestamp = 53;
        traffic_data[70].source_node = 12;
        traffic_data[70].dest_node = 15;
        traffic_data[70].packet_type = "CHI_READ";
        traffic_data[70].size_bytes = 64;
        traffic_data[71].timestamp = 53;
        traffic_data[71].source_node = 15;
        traffic_data[71].dest_node = 13;
        traffic_data[71].packet_type = "CHI_WRITE";
        traffic_data[71].size_bytes = 64;
        traffic_data[72].timestamp = 54;
        traffic_data[72].source_node = 7;
        traffic_data[72].dest_node = 15;
        traffic_data[72].packet_type = "AXI_WRITE";
        traffic_data[72].size_bytes = 64;
        traffic_data[73].timestamp = 55;
        traffic_data[73].source_node = 14;
        traffic_data[73].dest_node = 4;
        traffic_data[73].packet_type = "AXI_WRITE";
        traffic_data[73].size_bytes = 64;
        traffic_data[74].timestamp = 56;
        traffic_data[74].source_node = 2;
        traffic_data[74].dest_node = 4;
        traffic_data[74].packet_type = "AXI_READ";
        traffic_data[74].size_bytes = 64;
        traffic_data[75].timestamp = 56;
        traffic_data[75].source_node = 3;
        traffic_data[75].dest_node = 6;
        traffic_data[75].packet_type = "AXI_WRITE";
        traffic_data[75].size_bytes = 64;
        traffic_data[76].timestamp = 57;
        traffic_data[76].source_node = 10;
        traffic_data[76].dest_node = 4;
        traffic_data[76].packet_type = "AXI_READ";
        traffic_data[76].size_bytes = 64;
        traffic_data[77].timestamp = 57;
        traffic_data[77].source_node = 14;
        traffic_data[77].dest_node = 7;
        traffic_data[77].packet_type = "CHI_READ";
        traffic_data[77].size_bytes = 64;
        traffic_data[78].timestamp = 58;
        traffic_data[78].source_node = 3;
        traffic_data[78].dest_node = 13;
        traffic_data[78].packet_type = "CHI_READ";
        traffic_data[78].size_bytes = 64;
        traffic_data[79].timestamp = 58;
        traffic_data[79].source_node = 6;
        traffic_data[79].dest_node = 8;
        traffic_data[79].packet_type = "CHI_WRITE";
        traffic_data[79].size_bytes = 64;
        traffic_data[80].timestamp = 60;
        traffic_data[80].source_node = 9;
        traffic_data[80].dest_node = 1;
        traffic_data[80].packet_type = "AXI_READ";
        traffic_data[80].size_bytes = 64;
        traffic_data[81].timestamp = 60;
        traffic_data[81].source_node = 14;
        traffic_data[81].dest_node = 8;
        traffic_data[81].packet_type = "CHI_READ";
        traffic_data[81].size_bytes = 64;
        traffic_data[82].timestamp = 61;
        traffic_data[82].source_node = 5;
        traffic_data[82].dest_node = 4;
        traffic_data[82].packet_type = "CHI_READ";
        traffic_data[82].size_bytes = 64;
        traffic_data[83].timestamp = 62;
        traffic_data[83].source_node = 6;
        traffic_data[83].dest_node = 15;
        traffic_data[83].packet_type = "CHI_READ";
        traffic_data[83].size_bytes = 64;
        traffic_data[84].timestamp = 62;
        traffic_data[84].source_node = 7;
        traffic_data[84].dest_node = 4;
        traffic_data[84].packet_type = "CHI_READ";
        traffic_data[84].size_bytes = 64;
        traffic_data[85].timestamp = 62;
        traffic_data[85].source_node = 13;
        traffic_data[85].dest_node = 11;
        traffic_data[85].packet_type = "AXI_READ";
        traffic_data[85].size_bytes = 64;
        traffic_data[86].timestamp = 62;
        traffic_data[86].source_node = 14;
        traffic_data[86].dest_node = 8;
        traffic_data[86].packet_type = "AXI_WRITE";
        traffic_data[86].size_bytes = 64;
        traffic_data[87].timestamp = 63;
        traffic_data[87].source_node = 9;
        traffic_data[87].dest_node = 1;
        traffic_data[87].packet_type = "CHI_READ";
        traffic_data[87].size_bytes = 64;
        traffic_data[88].timestamp = 64;
        traffic_data[88].source_node = 8;
        traffic_data[88].dest_node = 3;
        traffic_data[88].packet_type = "CHI_READ";
        traffic_data[88].size_bytes = 64;
        traffic_data[89].timestamp = 65;
        traffic_data[89].source_node = 10;
        traffic_data[89].dest_node = 5;
        traffic_data[89].packet_type = "CHI_WRITE";
        traffic_data[89].size_bytes = 64;
        traffic_data[90].timestamp = 65;
        traffic_data[90].source_node = 15;
        traffic_data[90].dest_node = 5;
        traffic_data[90].packet_type = "AXI_WRITE";
        traffic_data[90].size_bytes = 64;
        traffic_data[91].timestamp = 66;
        traffic_data[91].source_node = 4;
        traffic_data[91].dest_node = 14;
        traffic_data[91].packet_type = "AXI_READ";
        traffic_data[91].size_bytes = 64;
        traffic_data[92].timestamp = 68;
        traffic_data[92].source_node = 8;
        traffic_data[92].dest_node = 7;
        traffic_data[92].packet_type = "CHI_READ";
        traffic_data[92].size_bytes = 64;
        traffic_data[93].timestamp = 68;
        traffic_data[93].source_node = 12;
        traffic_data[93].dest_node = 7;
        traffic_data[93].packet_type = "CHI_WRITE";
        traffic_data[93].size_bytes = 64;
        traffic_data[94].timestamp = 68;
        traffic_data[94].source_node = 13;
        traffic_data[94].dest_node = 5;
        traffic_data[94].packet_type = "CHI_READ";
        traffic_data[94].size_bytes = 64;
        traffic_data[95].timestamp = 68;
        traffic_data[95].source_node = 14;
        traffic_data[95].dest_node = 13;
        traffic_data[95].packet_type = "AXI_READ";
        traffic_data[95].size_bytes = 64;
        traffic_data[96].timestamp = 69;
        traffic_data[96].source_node = 11;
        traffic_data[96].dest_node = 1;
        traffic_data[96].packet_type = "CHI_READ";
        traffic_data[96].size_bytes = 64;
        traffic_data[97].timestamp = 69;
        traffic_data[97].source_node = 13;
        traffic_data[97].dest_node = 10;
        traffic_data[97].packet_type = "AXI_WRITE";
        traffic_data[97].size_bytes = 64;
        traffic_data[98].timestamp = 69;
        traffic_data[98].source_node = 14;
        traffic_data[98].dest_node = 11;
        traffic_data[98].packet_type = "CHI_WRITE";
        traffic_data[98].size_bytes = 64;
        traffic_data[99].timestamp = 70;
        traffic_data[99].source_node = 7;
        traffic_data[99].dest_node = 11;
        traffic_data[99].packet_type = "CHI_READ";
        traffic_data[99].size_bytes = 64;
        traffic_data[100].timestamp = 70;
        traffic_data[100].source_node = 8;
        traffic_data[100].dest_node = 1;
        traffic_data[100].packet_type = "CHI_WRITE";
        traffic_data[100].size_bytes = 64;
        traffic_data[101].timestamp = 72;
        traffic_data[101].source_node = 10;
        traffic_data[101].dest_node = 14;
        traffic_data[101].packet_type = "AXI_READ";
        traffic_data[101].size_bytes = 64;
        traffic_data[102].timestamp = 73;
        traffic_data[102].source_node = 9;
        traffic_data[102].dest_node = 5;
        traffic_data[102].packet_type = "AXI_WRITE";
        traffic_data[102].size_bytes = 64;
        traffic_data[103].timestamp = 74;
        traffic_data[103].source_node = 15;
        traffic_data[103].dest_node = 7;
        traffic_data[103].packet_type = "CHI_READ";
        traffic_data[103].size_bytes = 64;
        traffic_data[104].timestamp = 75;
        traffic_data[104].source_node = 14;
        traffic_data[104].dest_node = 0;
        traffic_data[104].packet_type = "CHI_WRITE";
        traffic_data[104].size_bytes = 64;
        traffic_data[105].timestamp = 76;
        traffic_data[105].source_node = 3;
        traffic_data[105].dest_node = 15;
        traffic_data[105].packet_type = "AXI_READ";
        traffic_data[105].size_bytes = 64;
        traffic_data[106].timestamp = 76;
        traffic_data[106].source_node = 14;
        traffic_data[106].dest_node = 1;
        traffic_data[106].packet_type = "AXI_READ";
        traffic_data[106].size_bytes = 64;
        traffic_data[107].timestamp = 77;
        traffic_data[107].source_node = 7;
        traffic_data[107].dest_node = 6;
        traffic_data[107].packet_type = "CHI_WRITE";
        traffic_data[107].size_bytes = 64;
        traffic_data[108].timestamp = 77;
        traffic_data[108].source_node = 8;
        traffic_data[108].dest_node = 14;
        traffic_data[108].packet_type = "CHI_WRITE";
        traffic_data[108].size_bytes = 64;
        traffic_data[109].timestamp = 77;
        traffic_data[109].source_node = 10;
        traffic_data[109].dest_node = 8;
        traffic_data[109].packet_type = "AXI_WRITE";
        traffic_data[109].size_bytes = 64;
        traffic_data[110].timestamp = 77;
        traffic_data[110].source_node = 13;
        traffic_data[110].dest_node = 5;
        traffic_data[110].packet_type = "AXI_WRITE";
        traffic_data[110].size_bytes = 64;
        traffic_data[111].timestamp = 78;
        traffic_data[111].source_node = 7;
        traffic_data[111].dest_node = 14;
        traffic_data[111].packet_type = "CHI_WRITE";
        traffic_data[111].size_bytes = 64;
        traffic_data[112].timestamp = 78;
        traffic_data[112].source_node = 8;
        traffic_data[112].dest_node = 6;
        traffic_data[112].packet_type = "CHI_READ";
        traffic_data[112].size_bytes = 64;
        traffic_data[113].timestamp = 78;
        traffic_data[113].source_node = 10;
        traffic_data[113].dest_node = 13;
        traffic_data[113].packet_type = "AXI_READ";
        traffic_data[113].size_bytes = 64;
        traffic_data[114].timestamp = 79;
        traffic_data[114].source_node = 1;
        traffic_data[114].dest_node = 9;
        traffic_data[114].packet_type = "CHI_READ";
        traffic_data[114].size_bytes = 64;
        traffic_data[115].timestamp = 79;
        traffic_data[115].source_node = 9;
        traffic_data[115].dest_node = 13;
        traffic_data[115].packet_type = "CHI_WRITE";
        traffic_data[115].size_bytes = 64;
        traffic_data[116].timestamp = 79;
        traffic_data[116].source_node = 10;
        traffic_data[116].dest_node = 3;
        traffic_data[116].packet_type = "AXI_READ";
        traffic_data[116].size_bytes = 64;
        traffic_data[117].timestamp = 80;
        traffic_data[117].source_node = 2;
        traffic_data[117].dest_node = 11;
        traffic_data[117].packet_type = "AXI_WRITE";
        traffic_data[117].size_bytes = 64;
        traffic_data[118].timestamp = 80;
        traffic_data[118].source_node = 5;
        traffic_data[118].dest_node = 11;
        traffic_data[118].packet_type = "CHI_READ";
        traffic_data[118].size_bytes = 64;
        traffic_data[119].timestamp = 81;
        traffic_data[119].source_node = 2;
        traffic_data[119].dest_node = 7;
        traffic_data[119].packet_type = "AXI_READ";
        traffic_data[119].size_bytes = 64;
        traffic_data[120].timestamp = 82;
        traffic_data[120].source_node = 5;
        traffic_data[120].dest_node = 11;
        traffic_data[120].packet_type = "CHI_WRITE";
        traffic_data[120].size_bytes = 64;
        traffic_data[121].timestamp = 82;
        traffic_data[121].source_node = 13;
        traffic_data[121].dest_node = 1;
        traffic_data[121].packet_type = "AXI_WRITE";
        traffic_data[121].size_bytes = 64;
        traffic_data[122].timestamp = 84;
        traffic_data[122].source_node = 13;
        traffic_data[122].dest_node = 10;
        traffic_data[122].packet_type = "CHI_READ";
        traffic_data[122].size_bytes = 64;
        traffic_data[123].timestamp = 86;
        traffic_data[123].source_node = 3;
        traffic_data[123].dest_node = 7;
        traffic_data[123].packet_type = "CHI_WRITE";
        traffic_data[123].size_bytes = 64;
        traffic_data[124].timestamp = 86;
        traffic_data[124].source_node = 7;
        traffic_data[124].dest_node = 5;
        traffic_data[124].packet_type = "AXI_READ";
        traffic_data[124].size_bytes = 64;
        traffic_data[125].timestamp = 87;
        traffic_data[125].source_node = 2;
        traffic_data[125].dest_node = 1;
        traffic_data[125].packet_type = "AXI_WRITE";
        traffic_data[125].size_bytes = 64;
        traffic_data[126].timestamp = 87;
        traffic_data[126].source_node = 10;
        traffic_data[126].dest_node = 3;
        traffic_data[126].packet_type = "CHI_READ";
        traffic_data[126].size_bytes = 64;
        traffic_data[127].timestamp = 88;
        traffic_data[127].source_node = 8;
        traffic_data[127].dest_node = 0;
        traffic_data[127].packet_type = "CHI_READ";
        traffic_data[127].size_bytes = 64;
        traffic_data[128].timestamp = 89;
        traffic_data[128].source_node = 5;
        traffic_data[128].dest_node = 0;
        traffic_data[128].packet_type = "AXI_WRITE";
        traffic_data[128].size_bytes = 64;
        traffic_data[129].timestamp = 90;
        traffic_data[129].source_node = 6;
        traffic_data[129].dest_node = 4;
        traffic_data[129].packet_type = "CHI_WRITE";
        traffic_data[129].size_bytes = 64;
        traffic_data[130].timestamp = 91;
        traffic_data[130].source_node = 4;
        traffic_data[130].dest_node = 7;
        traffic_data[130].packet_type = "CHI_WRITE";
        traffic_data[130].size_bytes = 64;
        traffic_data[131].timestamp = 91;
        traffic_data[131].source_node = 8;
        traffic_data[131].dest_node = 7;
        traffic_data[131].packet_type = "CHI_WRITE";
        traffic_data[131].size_bytes = 64;
        traffic_data[132].timestamp = 91;
        traffic_data[132].source_node = 10;
        traffic_data[132].dest_node = 1;
        traffic_data[132].packet_type = "CHI_WRITE";
        traffic_data[132].size_bytes = 64;
        traffic_data[133].timestamp = 91;
        traffic_data[133].source_node = 15;
        traffic_data[133].dest_node = 0;
        traffic_data[133].packet_type = "AXI_WRITE";
        traffic_data[133].size_bytes = 64;
        traffic_data[134].timestamp = 92;
        traffic_data[134].source_node = 9;
        traffic_data[134].dest_node = 5;
        traffic_data[134].packet_type = "CHI_READ";
        traffic_data[134].size_bytes = 64;
        traffic_data[135].timestamp = 92;
        traffic_data[135].source_node = 15;
        traffic_data[135].dest_node = 0;
        traffic_data[135].packet_type = "AXI_WRITE";
        traffic_data[135].size_bytes = 64;
        traffic_data[136].timestamp = 94;
        traffic_data[136].source_node = 1;
        traffic_data[136].dest_node = 6;
        traffic_data[136].packet_type = "AXI_READ";
        traffic_data[136].size_bytes = 64;
        traffic_data[137].timestamp = 94;
        traffic_data[137].source_node = 7;
        traffic_data[137].dest_node = 8;
        traffic_data[137].packet_type = "CHI_READ";
        traffic_data[137].size_bytes = 64;
        traffic_data[138].timestamp = 95;
        traffic_data[138].source_node = 4;
        traffic_data[138].dest_node = 12;
        traffic_data[138].packet_type = "AXI_READ";
        traffic_data[138].size_bytes = 64;
        traffic_data[139].timestamp = 98;
        traffic_data[139].source_node = 4;
        traffic_data[139].dest_node = 12;
        traffic_data[139].packet_type = "AXI_READ";
        traffic_data[139].size_bytes = 64;
        traffic_data[140].timestamp = 99;
        traffic_data[140].source_node = 4;
        traffic_data[140].dest_node = 7;
        traffic_data[140].packet_type = "CHI_READ";
        traffic_data[140].size_bytes = 64;
        traffic_data[141].timestamp = 99;
        traffic_data[141].source_node = 8;
        traffic_data[141].dest_node = 9;
        traffic_data[141].packet_type = "AXI_WRITE";
        traffic_data[141].size_bytes = 64;
        traffic_data[142].timestamp = 100;
        traffic_data[142].source_node = 2;
        traffic_data[142].dest_node = 10;
        traffic_data[142].packet_type = "AXI_WRITE";
        traffic_data[142].size_bytes = 64;
        traffic_data[143].timestamp = 101;
        traffic_data[143].source_node = 2;
        traffic_data[143].dest_node = 10;
        traffic_data[143].packet_type = "AXI_READ";
        traffic_data[143].size_bytes = 64;
        traffic_data[144].timestamp = 102;
        traffic_data[144].source_node = 1;
        traffic_data[144].dest_node = 6;
        traffic_data[144].packet_type = "CHI_READ";
        traffic_data[144].size_bytes = 64;
        traffic_data[145].timestamp = 102;
        traffic_data[145].source_node = 9;
        traffic_data[145].dest_node = 11;
        traffic_data[145].packet_type = "AXI_READ";
        traffic_data[145].size_bytes = 64;
        traffic_data[146].timestamp = 103;
        traffic_data[146].source_node = 4;
        traffic_data[146].dest_node = 11;
        traffic_data[146].packet_type = "CHI_READ";
        traffic_data[146].size_bytes = 64;
        traffic_data[147].timestamp = 103;
        traffic_data[147].source_node = 6;
        traffic_data[147].dest_node = 1;
        traffic_data[147].packet_type = "CHI_WRITE";
        traffic_data[147].size_bytes = 64;
        traffic_data[148].timestamp = 104;
        traffic_data[148].source_node = 15;
        traffic_data[148].dest_node = 7;
        traffic_data[148].packet_type = "CHI_READ";
        traffic_data[148].size_bytes = 64;
        traffic_data[149].timestamp = 105;
        traffic_data[149].source_node = 0;
        traffic_data[149].dest_node = 10;
        traffic_data[149].packet_type = "AXI_READ";
        traffic_data[149].size_bytes = 64;
        traffic_data[150].timestamp = 105;
        traffic_data[150].source_node = 1;
        traffic_data[150].dest_node = 9;
        traffic_data[150].packet_type = "AXI_WRITE";
        traffic_data[150].size_bytes = 64;
        traffic_data[151].timestamp = 105;
        traffic_data[151].source_node = 9;
        traffic_data[151].dest_node = 8;
        traffic_data[151].packet_type = "CHI_WRITE";
        traffic_data[151].size_bytes = 64;
        traffic_data[152].timestamp = 105;
        traffic_data[152].source_node = 14;
        traffic_data[152].dest_node = 7;
        traffic_data[152].packet_type = "CHI_READ";
        traffic_data[152].size_bytes = 64;
        traffic_data[153].timestamp = 106;
        traffic_data[153].source_node = 4;
        traffic_data[153].dest_node = 6;
        traffic_data[153].packet_type = "AXI_READ";
        traffic_data[153].size_bytes = 64;
        traffic_data[154].timestamp = 106;
        traffic_data[154].source_node = 6;
        traffic_data[154].dest_node = 15;
        traffic_data[154].packet_type = "AXI_READ";
        traffic_data[154].size_bytes = 64;
        traffic_data[155].timestamp = 107;
        traffic_data[155].source_node = 4;
        traffic_data[155].dest_node = 11;
        traffic_data[155].packet_type = "AXI_WRITE";
        traffic_data[155].size_bytes = 64;
        traffic_data[156].timestamp = 107;
        traffic_data[156].source_node = 12;
        traffic_data[156].dest_node = 0;
        traffic_data[156].packet_type = "CHI_READ";
        traffic_data[156].size_bytes = 64;
        traffic_data[157].timestamp = 108;
        traffic_data[157].source_node = 7;
        traffic_data[157].dest_node = 11;
        traffic_data[157].packet_type = "CHI_WRITE";
        traffic_data[157].size_bytes = 64;
        traffic_data[158].timestamp = 108;
        traffic_data[158].source_node = 12;
        traffic_data[158].dest_node = 9;
        traffic_data[158].packet_type = "AXI_READ";
        traffic_data[158].size_bytes = 64;
        traffic_data[159].timestamp = 109;
        traffic_data[159].source_node = 1;
        traffic_data[159].dest_node = 8;
        traffic_data[159].packet_type = "AXI_WRITE";
        traffic_data[159].size_bytes = 64;
        traffic_data[160].timestamp = 110;
        traffic_data[160].source_node = 9;
        traffic_data[160].dest_node = 5;
        traffic_data[160].packet_type = "CHI_WRITE";
        traffic_data[160].size_bytes = 64;
        traffic_data[161].timestamp = 111;
        traffic_data[161].source_node = 15;
        traffic_data[161].dest_node = 11;
        traffic_data[161].packet_type = "AXI_WRITE";
        traffic_data[161].size_bytes = 64;
        traffic_data[162].timestamp = 112;
        traffic_data[162].source_node = 0;
        traffic_data[162].dest_node = 7;
        traffic_data[162].packet_type = "AXI_READ";
        traffic_data[162].size_bytes = 64;
        traffic_data[163].timestamp = 112;
        traffic_data[163].source_node = 10;
        traffic_data[163].dest_node = 15;
        traffic_data[163].packet_type = "AXI_WRITE";
        traffic_data[163].size_bytes = 64;
        traffic_data[164].timestamp = 113;
        traffic_data[164].source_node = 11;
        traffic_data[164].dest_node = 12;
        traffic_data[164].packet_type = "CHI_WRITE";
        traffic_data[164].size_bytes = 64;
        traffic_data[165].timestamp = 114;
        traffic_data[165].source_node = 0;
        traffic_data[165].dest_node = 14;
        traffic_data[165].packet_type = "AXI_WRITE";
        traffic_data[165].size_bytes = 64;
        traffic_data[166].timestamp = 114;
        traffic_data[166].source_node = 2;
        traffic_data[166].dest_node = 9;
        traffic_data[166].packet_type = "CHI_WRITE";
        traffic_data[166].size_bytes = 64;
        traffic_data[167].timestamp = 115;
        traffic_data[167].source_node = 10;
        traffic_data[167].dest_node = 14;
        traffic_data[167].packet_type = "AXI_READ";
        traffic_data[167].size_bytes = 64;
        traffic_data[168].timestamp = 116;
        traffic_data[168].source_node = 0;
        traffic_data[168].dest_node = 9;
        traffic_data[168].packet_type = "CHI_WRITE";
        traffic_data[168].size_bytes = 64;
        traffic_data[169].timestamp = 116;
        traffic_data[169].source_node = 7;
        traffic_data[169].dest_node = 9;
        traffic_data[169].packet_type = "CHI_WRITE";
        traffic_data[169].size_bytes = 64;
        traffic_data[170].timestamp = 116;
        traffic_data[170].source_node = 8;
        traffic_data[170].dest_node = 9;
        traffic_data[170].packet_type = "CHI_READ";
        traffic_data[170].size_bytes = 64;
        traffic_data[171].timestamp = 117;
        traffic_data[171].source_node = 7;
        traffic_data[171].dest_node = 6;
        traffic_data[171].packet_type = "CHI_WRITE";
        traffic_data[171].size_bytes = 64;
        traffic_data[172].timestamp = 118;
        traffic_data[172].source_node = 0;
        traffic_data[172].dest_node = 7;
        traffic_data[172].packet_type = "CHI_WRITE";
        traffic_data[172].size_bytes = 64;
        traffic_data[173].timestamp = 118;
        traffic_data[173].source_node = 2;
        traffic_data[173].dest_node = 0;
        traffic_data[173].packet_type = "AXI_WRITE";
        traffic_data[173].size_bytes = 64;
        traffic_data[174].timestamp = 118;
        traffic_data[174].source_node = 3;
        traffic_data[174].dest_node = 14;
        traffic_data[174].packet_type = "CHI_WRITE";
        traffic_data[174].size_bytes = 64;
        traffic_data[175].timestamp = 119;
        traffic_data[175].source_node = 6;
        traffic_data[175].dest_node = 3;
        traffic_data[175].packet_type = "AXI_WRITE";
        traffic_data[175].size_bytes = 64;
        traffic_data[176].timestamp = 119;
        traffic_data[176].source_node = 10;
        traffic_data[176].dest_node = 2;
        traffic_data[176].packet_type = "AXI_WRITE";
        traffic_data[176].size_bytes = 64;
        traffic_data[177].timestamp = 120;
        traffic_data[177].source_node = 3;
        traffic_data[177].dest_node = 12;
        traffic_data[177].packet_type = "CHI_READ";
        traffic_data[177].size_bytes = 64;
        traffic_data[178].timestamp = 120;
        traffic_data[178].source_node = 4;
        traffic_data[178].dest_node = 7;
        traffic_data[178].packet_type = "AXI_WRITE";
        traffic_data[178].size_bytes = 64;
        traffic_data[179].timestamp = 120;
        traffic_data[179].source_node = 11;
        traffic_data[179].dest_node = 4;
        traffic_data[179].packet_type = "CHI_WRITE";
        traffic_data[179].size_bytes = 64;
        traffic_data[180].timestamp = 121;
        traffic_data[180].source_node = 2;
        traffic_data[180].dest_node = 10;
        traffic_data[180].packet_type = "CHI_READ";
        traffic_data[180].size_bytes = 64;
        traffic_data[181].timestamp = 121;
        traffic_data[181].source_node = 5;
        traffic_data[181].dest_node = 2;
        traffic_data[181].packet_type = "CHI_WRITE";
        traffic_data[181].size_bytes = 64;
        traffic_data[182].timestamp = 121;
        traffic_data[182].source_node = 11;
        traffic_data[182].dest_node = 4;
        traffic_data[182].packet_type = "CHI_WRITE";
        traffic_data[182].size_bytes = 64;
        traffic_data[183].timestamp = 122;
        traffic_data[183].source_node = 3;
        traffic_data[183].dest_node = 6;
        traffic_data[183].packet_type = "AXI_READ";
        traffic_data[183].size_bytes = 64;
        traffic_data[184].timestamp = 122;
        traffic_data[184].source_node = 7;
        traffic_data[184].dest_node = 6;
        traffic_data[184].packet_type = "CHI_WRITE";
        traffic_data[184].size_bytes = 64;
        traffic_data[185].timestamp = 123;
        traffic_data[185].source_node = 14;
        traffic_data[185].dest_node = 6;
        traffic_data[185].packet_type = "CHI_READ";
        traffic_data[185].size_bytes = 64;
        traffic_data[186].timestamp = 125;
        traffic_data[186].source_node = 11;
        traffic_data[186].dest_node = 12;
        traffic_data[186].packet_type = "CHI_WRITE";
        traffic_data[186].size_bytes = 64;
        traffic_data[187].timestamp = 126;
        traffic_data[187].source_node = 0;
        traffic_data[187].dest_node = 14;
        traffic_data[187].packet_type = "CHI_WRITE";
        traffic_data[187].size_bytes = 64;
        traffic_data[188].timestamp = 126;
        traffic_data[188].source_node = 15;
        traffic_data[188].dest_node = 5;
        traffic_data[188].packet_type = "AXI_READ";
        traffic_data[188].size_bytes = 64;
        traffic_data[189].timestamp = 127;
        traffic_data[189].source_node = 12;
        traffic_data[189].dest_node = 3;
        traffic_data[189].packet_type = "AXI_WRITE";
        traffic_data[189].size_bytes = 64;
        traffic_data[190].timestamp = 128;
        traffic_data[190].source_node = 3;
        traffic_data[190].dest_node = 1;
        traffic_data[190].packet_type = "CHI_READ";
        traffic_data[190].size_bytes = 64;
        traffic_data[191].timestamp = 130;
        traffic_data[191].source_node = 3;
        traffic_data[191].dest_node = 10;
        traffic_data[191].packet_type = "AXI_WRITE";
        traffic_data[191].size_bytes = 64;
        traffic_data[192].timestamp = 130;
        traffic_data[192].source_node = 6;
        traffic_data[192].dest_node = 3;
        traffic_data[192].packet_type = "AXI_WRITE";
        traffic_data[192].size_bytes = 64;
        traffic_data[193].timestamp = 134;
        traffic_data[193].source_node = 1;
        traffic_data[193].dest_node = 4;
        traffic_data[193].packet_type = "CHI_READ";
        traffic_data[193].size_bytes = 64;
        traffic_data[194].timestamp = 134;
        traffic_data[194].source_node = 13;
        traffic_data[194].dest_node = 11;
        traffic_data[194].packet_type = "CHI_WRITE";
        traffic_data[194].size_bytes = 64;
        traffic_data[195].timestamp = 136;
        traffic_data[195].source_node = 5;
        traffic_data[195].dest_node = 6;
        traffic_data[195].packet_type = "CHI_READ";
        traffic_data[195].size_bytes = 64;
        traffic_data[196].timestamp = 137;
        traffic_data[196].source_node = 2;
        traffic_data[196].dest_node = 5;
        traffic_data[196].packet_type = "AXI_WRITE";
        traffic_data[196].size_bytes = 64;
        traffic_data[197].timestamp = 137;
        traffic_data[197].source_node = 14;
        traffic_data[197].dest_node = 12;
        traffic_data[197].packet_type = "AXI_READ";
        traffic_data[197].size_bytes = 64;
        traffic_data[198].timestamp = 138;
        traffic_data[198].source_node = 8;
        traffic_data[198].dest_node = 7;
        traffic_data[198].packet_type = "CHI_READ";
        traffic_data[198].size_bytes = 64;
        traffic_data[199].timestamp = 139;
        traffic_data[199].source_node = 7;
        traffic_data[199].dest_node = 11;
        traffic_data[199].packet_type = "CHI_WRITE";
        traffic_data[199].size_bytes = 64;
        traffic_data[200].timestamp = 139;
        traffic_data[200].source_node = 8;
        traffic_data[200].dest_node = 15;
        traffic_data[200].packet_type = "AXI_WRITE";
        traffic_data[200].size_bytes = 64;
        traffic_data[201].timestamp = 139;
        traffic_data[201].source_node = 10;
        traffic_data[201].dest_node = 6;
        traffic_data[201].packet_type = "AXI_WRITE";
        traffic_data[201].size_bytes = 64;
        traffic_data[202].timestamp = 140;
        traffic_data[202].source_node = 1;
        traffic_data[202].dest_node = 6;
        traffic_data[202].packet_type = "CHI_READ";
        traffic_data[202].size_bytes = 64;
        traffic_data[203].timestamp = 140;
        traffic_data[203].source_node = 2;
        traffic_data[203].dest_node = 11;
        traffic_data[203].packet_type = "AXI_WRITE";
        traffic_data[203].size_bytes = 64;
        traffic_data[204].timestamp = 140;
        traffic_data[204].source_node = 3;
        traffic_data[204].dest_node = 11;
        traffic_data[204].packet_type = "CHI_READ";
        traffic_data[204].size_bytes = 64;
        traffic_data[205].timestamp = 140;
        traffic_data[205].source_node = 7;
        traffic_data[205].dest_node = 1;
        traffic_data[205].packet_type = "AXI_READ";
        traffic_data[205].size_bytes = 64;
        traffic_data[206].timestamp = 140;
        traffic_data[206].source_node = 9;
        traffic_data[206].dest_node = 10;
        traffic_data[206].packet_type = "AXI_WRITE";
        traffic_data[206].size_bytes = 64;
        traffic_data[207].timestamp = 140;
        traffic_data[207].source_node = 12;
        traffic_data[207].dest_node = 5;
        traffic_data[207].packet_type = "AXI_READ";
        traffic_data[207].size_bytes = 64;
        traffic_data[208].timestamp = 141;
        traffic_data[208].source_node = 0;
        traffic_data[208].dest_node = 7;
        traffic_data[208].packet_type = "AXI_READ";
        traffic_data[208].size_bytes = 64;
        traffic_data[209].timestamp = 141;
        traffic_data[209].source_node = 12;
        traffic_data[209].dest_node = 10;
        traffic_data[209].packet_type = "AXI_WRITE";
        traffic_data[209].size_bytes = 64;
        traffic_data[210].timestamp = 142;
        traffic_data[210].source_node = 4;
        traffic_data[210].dest_node = 1;
        traffic_data[210].packet_type = "AXI_WRITE";
        traffic_data[210].size_bytes = 64;
        traffic_data[211].timestamp = 142;
        traffic_data[211].source_node = 12;
        traffic_data[211].dest_node = 8;
        traffic_data[211].packet_type = "CHI_READ";
        traffic_data[211].size_bytes = 64;
        traffic_data[212].timestamp = 143;
        traffic_data[212].source_node = 6;
        traffic_data[212].dest_node = 15;
        traffic_data[212].packet_type = "AXI_WRITE";
        traffic_data[212].size_bytes = 64;
        traffic_data[213].timestamp = 144;
        traffic_data[213].source_node = 7;
        traffic_data[213].dest_node = 1;
        traffic_data[213].packet_type = "AXI_READ";
        traffic_data[213].size_bytes = 64;
        traffic_data[214].timestamp = 144;
        traffic_data[214].source_node = 9;
        traffic_data[214].dest_node = 0;
        traffic_data[214].packet_type = "CHI_WRITE";
        traffic_data[214].size_bytes = 64;
        traffic_data[215].timestamp = 144;
        traffic_data[215].source_node = 15;
        traffic_data[215].dest_node = 8;
        traffic_data[215].packet_type = "AXI_WRITE";
        traffic_data[215].size_bytes = 64;
        traffic_data[216].timestamp = 145;
        traffic_data[216].source_node = 10;
        traffic_data[216].dest_node = 12;
        traffic_data[216].packet_type = "CHI_WRITE";
        traffic_data[216].size_bytes = 64;
        traffic_data[217].timestamp = 145;
        traffic_data[217].source_node = 13;
        traffic_data[217].dest_node = 1;
        traffic_data[217].packet_type = "CHI_WRITE";
        traffic_data[217].size_bytes = 64;
        traffic_data[218].timestamp = 146;
        traffic_data[218].source_node = 0;
        traffic_data[218].dest_node = 11;
        traffic_data[218].packet_type = "AXI_WRITE";
        traffic_data[218].size_bytes = 64;
        traffic_data[219].timestamp = 146;
        traffic_data[219].source_node = 15;
        traffic_data[219].dest_node = 12;
        traffic_data[219].packet_type = "CHI_WRITE";
        traffic_data[219].size_bytes = 64;
        traffic_data[220].timestamp = 147;
        traffic_data[220].source_node = 1;
        traffic_data[220].dest_node = 12;
        traffic_data[220].packet_type = "AXI_READ";
        traffic_data[220].size_bytes = 64;
        traffic_data[221].timestamp = 147;
        traffic_data[221].source_node = 4;
        traffic_data[221].dest_node = 14;
        traffic_data[221].packet_type = "AXI_WRITE";
        traffic_data[221].size_bytes = 64;
        traffic_data[222].timestamp = 147;
        traffic_data[222].source_node = 12;
        traffic_data[222].dest_node = 14;
        traffic_data[222].packet_type = "AXI_READ";
        traffic_data[222].size_bytes = 64;
        traffic_data[223].timestamp = 148;
        traffic_data[223].source_node = 11;
        traffic_data[223].dest_node = 5;
        traffic_data[223].packet_type = "AXI_READ";
        traffic_data[223].size_bytes = 64;
        traffic_data[224].timestamp = 149;
        traffic_data[224].source_node = 2;
        traffic_data[224].dest_node = 8;
        traffic_data[224].packet_type = "CHI_READ";
        traffic_data[224].size_bytes = 64;
        traffic_data[225].timestamp = 149;
        traffic_data[225].source_node = 5;
        traffic_data[225].dest_node = 8;
        traffic_data[225].packet_type = "AXI_READ";
        traffic_data[225].size_bytes = 64;
        traffic_data[226].timestamp = 150;
        traffic_data[226].source_node = 4;
        traffic_data[226].dest_node = 9;
        traffic_data[226].packet_type = "CHI_READ";
        traffic_data[226].size_bytes = 64;
        traffic_data[227].timestamp = 150;
        traffic_data[227].source_node = 7;
        traffic_data[227].dest_node = 5;
        traffic_data[227].packet_type = "AXI_READ";
        traffic_data[227].size_bytes = 64;
        traffic_data[228].timestamp = 151;
        traffic_data[228].source_node = 3;
        traffic_data[228].dest_node = 4;
        traffic_data[228].packet_type = "CHI_WRITE";
        traffic_data[228].size_bytes = 64;
        traffic_data[229].timestamp = 151;
        traffic_data[229].source_node = 7;
        traffic_data[229].dest_node = 1;
        traffic_data[229].packet_type = "AXI_WRITE";
        traffic_data[229].size_bytes = 64;
        traffic_data[230].timestamp = 151;
        traffic_data[230].source_node = 11;
        traffic_data[230].dest_node = 10;
        traffic_data[230].packet_type = "AXI_WRITE";
        traffic_data[230].size_bytes = 64;
        traffic_data[231].timestamp = 152;
        traffic_data[231].source_node = 4;
        traffic_data[231].dest_node = 3;
        traffic_data[231].packet_type = "AXI_WRITE";
        traffic_data[231].size_bytes = 64;
        traffic_data[232].timestamp = 153;
        traffic_data[232].source_node = 5;
        traffic_data[232].dest_node = 14;
        traffic_data[232].packet_type = "CHI_READ";
        traffic_data[232].size_bytes = 64;
        traffic_data[233].timestamp = 153;
        traffic_data[233].source_node = 10;
        traffic_data[233].dest_node = 4;
        traffic_data[233].packet_type = "CHI_READ";
        traffic_data[233].size_bytes = 64;
        traffic_data[234].timestamp = 154;
        traffic_data[234].source_node = 1;
        traffic_data[234].dest_node = 2;
        traffic_data[234].packet_type = "AXI_WRITE";
        traffic_data[234].size_bytes = 64;
        traffic_data[235].timestamp = 154;
        traffic_data[235].source_node = 3;
        traffic_data[235].dest_node = 13;
        traffic_data[235].packet_type = "AXI_WRITE";
        traffic_data[235].size_bytes = 64;
        traffic_data[236].timestamp = 154;
        traffic_data[236].source_node = 12;
        traffic_data[236].dest_node = 1;
        traffic_data[236].packet_type = "AXI_WRITE";
        traffic_data[236].size_bytes = 64;
        traffic_data[237].timestamp = 155;
        traffic_data[237].source_node = 3;
        traffic_data[237].dest_node = 8;
        traffic_data[237].packet_type = "AXI_READ";
        traffic_data[237].size_bytes = 64;
        traffic_data[238].timestamp = 155;
        traffic_data[238].source_node = 8;
        traffic_data[238].dest_node = 11;
        traffic_data[238].packet_type = "CHI_WRITE";
        traffic_data[238].size_bytes = 64;
        traffic_data[239].timestamp = 155;
        traffic_data[239].source_node = 14;
        traffic_data[239].dest_node = 9;
        traffic_data[239].packet_type = "AXI_WRITE";
        traffic_data[239].size_bytes = 64;
        traffic_data[240].timestamp = 156;
        traffic_data[240].source_node = 3;
        traffic_data[240].dest_node = 7;
        traffic_data[240].packet_type = "AXI_WRITE";
        traffic_data[240].size_bytes = 64;
        traffic_data[241].timestamp = 156;
        traffic_data[241].source_node = 10;
        traffic_data[241].dest_node = 6;
        traffic_data[241].packet_type = "CHI_READ";
        traffic_data[241].size_bytes = 64;
        traffic_data[242].timestamp = 157;
        traffic_data[242].source_node = 1;
        traffic_data[242].dest_node = 10;
        traffic_data[242].packet_type = "AXI_WRITE";
        traffic_data[242].size_bytes = 64;
        traffic_data[243].timestamp = 157;
        traffic_data[243].source_node = 2;
        traffic_data[243].dest_node = 13;
        traffic_data[243].packet_type = "CHI_READ";
        traffic_data[243].size_bytes = 64;
        traffic_data[244].timestamp = 157;
        traffic_data[244].source_node = 3;
        traffic_data[244].dest_node = 8;
        traffic_data[244].packet_type = "CHI_READ";
        traffic_data[244].size_bytes = 64;
        traffic_data[245].timestamp = 157;
        traffic_data[245].source_node = 12;
        traffic_data[245].dest_node = 3;
        traffic_data[245].packet_type = "CHI_WRITE";
        traffic_data[245].size_bytes = 64;
        traffic_data[246].timestamp = 158;
        traffic_data[246].source_node = 5;
        traffic_data[246].dest_node = 12;
        traffic_data[246].packet_type = "CHI_READ";
        traffic_data[246].size_bytes = 64;
        traffic_data[247].timestamp = 158;
        traffic_data[247].source_node = 15;
        traffic_data[247].dest_node = 3;
        traffic_data[247].packet_type = "AXI_WRITE";
        traffic_data[247].size_bytes = 64;
        traffic_data[248].timestamp = 159;
        traffic_data[248].source_node = 0;
        traffic_data[248].dest_node = 8;
        traffic_data[248].packet_type = "AXI_READ";
        traffic_data[248].size_bytes = 64;
        traffic_data[249].timestamp = 159;
        traffic_data[249].source_node = 8;
        traffic_data[249].dest_node = 2;
        traffic_data[249].packet_type = "AXI_WRITE";
        traffic_data[249].size_bytes = 64;
        traffic_data[250].timestamp = 161;
        traffic_data[250].source_node = 9;
        traffic_data[250].dest_node = 10;
        traffic_data[250].packet_type = "CHI_READ";
        traffic_data[250].size_bytes = 64;
        traffic_data[251].timestamp = 162;
        traffic_data[251].source_node = 5;
        traffic_data[251].dest_node = 12;
        traffic_data[251].packet_type = "CHI_READ";
        traffic_data[251].size_bytes = 64;
        traffic_data[252].timestamp = 162;
        traffic_data[252].source_node = 9;
        traffic_data[252].dest_node = 4;
        traffic_data[252].packet_type = "AXI_READ";
        traffic_data[252].size_bytes = 64;
        traffic_data[253].timestamp = 162;
        traffic_data[253].source_node = 11;
        traffic_data[253].dest_node = 7;
        traffic_data[253].packet_type = "CHI_WRITE";
        traffic_data[253].size_bytes = 64;
        traffic_data[254].timestamp = 163;
        traffic_data[254].source_node = 7;
        traffic_data[254].dest_node = 14;
        traffic_data[254].packet_type = "AXI_READ";
        traffic_data[254].size_bytes = 64;
        traffic_data[255].timestamp = 163;
        traffic_data[255].source_node = 11;
        traffic_data[255].dest_node = 2;
        traffic_data[255].packet_type = "CHI_WRITE";
        traffic_data[255].size_bytes = 64;
        traffic_data[256].timestamp = 163;
        traffic_data[256].source_node = 13;
        traffic_data[256].dest_node = 15;
        traffic_data[256].packet_type = "AXI_READ";
        traffic_data[256].size_bytes = 64;
        traffic_data[257].timestamp = 164;
        traffic_data[257].source_node = 6;
        traffic_data[257].dest_node = 5;
        traffic_data[257].packet_type = "AXI_WRITE";
        traffic_data[257].size_bytes = 64;
        traffic_data[258].timestamp = 164;
        traffic_data[258].source_node = 14;
        traffic_data[258].dest_node = 6;
        traffic_data[258].packet_type = "CHI_WRITE";
        traffic_data[258].size_bytes = 64;
        traffic_data[259].timestamp = 165;
        traffic_data[259].source_node = 6;
        traffic_data[259].dest_node = 2;
        traffic_data[259].packet_type = "CHI_READ";
        traffic_data[259].size_bytes = 64;
        traffic_data[260].timestamp = 166;
        traffic_data[260].source_node = 3;
        traffic_data[260].dest_node = 8;
        traffic_data[260].packet_type = "CHI_WRITE";
        traffic_data[260].size_bytes = 64;
        traffic_data[261].timestamp = 166;
        traffic_data[261].source_node = 9;
        traffic_data[261].dest_node = 11;
        traffic_data[261].packet_type = "CHI_READ";
        traffic_data[261].size_bytes = 64;
        traffic_data[262].timestamp = 166;
        traffic_data[262].source_node = 14;
        traffic_data[262].dest_node = 6;
        traffic_data[262].packet_type = "CHI_WRITE";
        traffic_data[262].size_bytes = 64;
        traffic_data[263].timestamp = 167;
        traffic_data[263].source_node = 7;
        traffic_data[263].dest_node = 10;
        traffic_data[263].packet_type = "AXI_WRITE";
        traffic_data[263].size_bytes = 64;
        traffic_data[264].timestamp = 168;
        traffic_data[264].source_node = 8;
        traffic_data[264].dest_node = 6;
        traffic_data[264].packet_type = "CHI_WRITE";
        traffic_data[264].size_bytes = 64;
        traffic_data[265].timestamp = 168;
        traffic_data[265].source_node = 13;
        traffic_data[265].dest_node = 11;
        traffic_data[265].packet_type = "CHI_WRITE";
        traffic_data[265].size_bytes = 64;
        traffic_data[266].timestamp = 170;
        traffic_data[266].source_node = 6;
        traffic_data[266].dest_node = 8;
        traffic_data[266].packet_type = "CHI_READ";
        traffic_data[266].size_bytes = 64;
        traffic_data[267].timestamp = 170;
        traffic_data[267].source_node = 8;
        traffic_data[267].dest_node = 14;
        traffic_data[267].packet_type = "CHI_READ";
        traffic_data[267].size_bytes = 64;
        traffic_data[268].timestamp = 171;
        traffic_data[268].source_node = 5;
        traffic_data[268].dest_node = 8;
        traffic_data[268].packet_type = "AXI_WRITE";
        traffic_data[268].size_bytes = 64;
        traffic_data[269].timestamp = 171;
        traffic_data[269].source_node = 11;
        traffic_data[269].dest_node = 13;
        traffic_data[269].packet_type = "AXI_WRITE";
        traffic_data[269].size_bytes = 64;
        traffic_data[270].timestamp = 171;
        traffic_data[270].source_node = 12;
        traffic_data[270].dest_node = 11;
        traffic_data[270].packet_type = "CHI_WRITE";
        traffic_data[270].size_bytes = 64;
        traffic_data[271].timestamp = 172;
        traffic_data[271].source_node = 0;
        traffic_data[271].dest_node = 4;
        traffic_data[271].packet_type = "AXI_WRITE";
        traffic_data[271].size_bytes = 64;
        traffic_data[272].timestamp = 172;
        traffic_data[272].source_node = 11;
        traffic_data[272].dest_node = 5;
        traffic_data[272].packet_type = "CHI_WRITE";
        traffic_data[272].size_bytes = 64;
        traffic_data[273].timestamp = 173;
        traffic_data[273].source_node = 15;
        traffic_data[273].dest_node = 12;
        traffic_data[273].packet_type = "AXI_READ";
        traffic_data[273].size_bytes = 64;
        traffic_data[274].timestamp = 175;
        traffic_data[274].source_node = 2;
        traffic_data[274].dest_node = 11;
        traffic_data[274].packet_type = "CHI_READ";
        traffic_data[274].size_bytes = 64;
        traffic_data[275].timestamp = 176;
        traffic_data[275].source_node = 2;
        traffic_data[275].dest_node = 14;
        traffic_data[275].packet_type = "CHI_WRITE";
        traffic_data[275].size_bytes = 64;
        traffic_data[276].timestamp = 176;
        traffic_data[276].source_node = 11;
        traffic_data[276].dest_node = 12;
        traffic_data[276].packet_type = "AXI_WRITE";
        traffic_data[276].size_bytes = 64;
        traffic_data[277].timestamp = 178;
        traffic_data[277].source_node = 9;
        traffic_data[277].dest_node = 11;
        traffic_data[277].packet_type = "AXI_READ";
        traffic_data[277].size_bytes = 64;
        traffic_data[278].timestamp = 179;
        traffic_data[278].source_node = 10;
        traffic_data[278].dest_node = 5;
        traffic_data[278].packet_type = "AXI_WRITE";
        traffic_data[278].size_bytes = 64;
        traffic_data[279].timestamp = 179;
        traffic_data[279].source_node = 12;
        traffic_data[279].dest_node = 7;
        traffic_data[279].packet_type = "CHI_READ";
        traffic_data[279].size_bytes = 64;
        traffic_data[280].timestamp = 180;
        traffic_data[280].source_node = 8;
        traffic_data[280].dest_node = 9;
        traffic_data[280].packet_type = "AXI_WRITE";
        traffic_data[280].size_bytes = 64;
        traffic_data[281].timestamp = 180;
        traffic_data[281].source_node = 14;
        traffic_data[281].dest_node = 0;
        traffic_data[281].packet_type = "AXI_WRITE";
        traffic_data[281].size_bytes = 64;
        traffic_data[282].timestamp = 181;
        traffic_data[282].source_node = 5;
        traffic_data[282].dest_node = 0;
        traffic_data[282].packet_type = "CHI_READ";
        traffic_data[282].size_bytes = 64;
        traffic_data[283].timestamp = 182;
        traffic_data[283].source_node = 3;
        traffic_data[283].dest_node = 4;
        traffic_data[283].packet_type = "AXI_WRITE";
        traffic_data[283].size_bytes = 64;
        traffic_data[284].timestamp = 182;
        traffic_data[284].source_node = 5;
        traffic_data[284].dest_node = 9;
        traffic_data[284].packet_type = "AXI_WRITE";
        traffic_data[284].size_bytes = 64;
        traffic_data[285].timestamp = 182;
        traffic_data[285].source_node = 14;
        traffic_data[285].dest_node = 1;
        traffic_data[285].packet_type = "AXI_READ";
        traffic_data[285].size_bytes = 64;
        traffic_data[286].timestamp = 182;
        traffic_data[286].source_node = 15;
        traffic_data[286].dest_node = 1;
        traffic_data[286].packet_type = "CHI_WRITE";
        traffic_data[286].size_bytes = 64;
        traffic_data[287].timestamp = 183;
        traffic_data[287].source_node = 6;
        traffic_data[287].dest_node = 7;
        traffic_data[287].packet_type = "AXI_READ";
        traffic_data[287].size_bytes = 64;
        traffic_data[288].timestamp = 184;
        traffic_data[288].source_node = 8;
        traffic_data[288].dest_node = 7;
        traffic_data[288].packet_type = "AXI_WRITE";
        traffic_data[288].size_bytes = 64;
        traffic_data[289].timestamp = 184;
        traffic_data[289].source_node = 12;
        traffic_data[289].dest_node = 1;
        traffic_data[289].packet_type = "AXI_READ";
        traffic_data[289].size_bytes = 64;
        traffic_data[290].timestamp = 185;
        traffic_data[290].source_node = 0;
        traffic_data[290].dest_node = 9;
        traffic_data[290].packet_type = "AXI_READ";
        traffic_data[290].size_bytes = 64;
        traffic_data[291].timestamp = 185;
        traffic_data[291].source_node = 8;
        traffic_data[291].dest_node = 2;
        traffic_data[291].packet_type = "AXI_READ";
        traffic_data[291].size_bytes = 64;
        traffic_data[292].timestamp = 186;
        traffic_data[292].source_node = 0;
        traffic_data[292].dest_node = 3;
        traffic_data[292].packet_type = "AXI_WRITE";
        traffic_data[292].size_bytes = 64;
        traffic_data[293].timestamp = 188;
        traffic_data[293].source_node = 5;
        traffic_data[293].dest_node = 11;
        traffic_data[293].packet_type = "CHI_READ";
        traffic_data[293].size_bytes = 64;
        traffic_data[294].timestamp = 188;
        traffic_data[294].source_node = 6;
        traffic_data[294].dest_node = 14;
        traffic_data[294].packet_type = "AXI_WRITE";
        traffic_data[294].size_bytes = 64;
        traffic_data[295].timestamp = 188;
        traffic_data[295].source_node = 12;
        traffic_data[295].dest_node = 10;
        traffic_data[295].packet_type = "AXI_WRITE";
        traffic_data[295].size_bytes = 64;
        traffic_data[296].timestamp = 189;
        traffic_data[296].source_node = 4;
        traffic_data[296].dest_node = 15;
        traffic_data[296].packet_type = "AXI_WRITE";
        traffic_data[296].size_bytes = 64;
        traffic_data[297].timestamp = 190;
        traffic_data[297].source_node = 1;
        traffic_data[297].dest_node = 8;
        traffic_data[297].packet_type = "CHI_WRITE";
        traffic_data[297].size_bytes = 64;
        traffic_data[298].timestamp = 190;
        traffic_data[298].source_node = 2;
        traffic_data[298].dest_node = 8;
        traffic_data[298].packet_type = "CHI_WRITE";
        traffic_data[298].size_bytes = 64;
        traffic_data[299].timestamp = 190;
        traffic_data[299].source_node = 6;
        traffic_data[299].dest_node = 7;
        traffic_data[299].packet_type = "CHI_WRITE";
        traffic_data[299].size_bytes = 64;
        traffic_data[300].timestamp = 190;
        traffic_data[300].source_node = 7;
        traffic_data[300].dest_node = 9;
        traffic_data[300].packet_type = "AXI_READ";
        traffic_data[300].size_bytes = 64;
        traffic_data[301].timestamp = 191;
        traffic_data[301].source_node = 10;
        traffic_data[301].dest_node = 11;
        traffic_data[301].packet_type = "AXI_WRITE";
        traffic_data[301].size_bytes = 64;
        traffic_data[302].timestamp = 191;
        traffic_data[302].source_node = 11;
        traffic_data[302].dest_node = 5;
        traffic_data[302].packet_type = "CHI_READ";
        traffic_data[302].size_bytes = 64;
        traffic_data[303].timestamp = 192;
        traffic_data[303].source_node = 13;
        traffic_data[303].dest_node = 10;
        traffic_data[303].packet_type = "AXI_READ";
        traffic_data[303].size_bytes = 64;
        traffic_data[304].timestamp = 193;
        traffic_data[304].source_node = 5;
        traffic_data[304].dest_node = 15;
        traffic_data[304].packet_type = "CHI_WRITE";
        traffic_data[304].size_bytes = 64;
        traffic_data[305].timestamp = 196;
        traffic_data[305].source_node = 11;
        traffic_data[305].dest_node = 2;
        traffic_data[305].packet_type = "AXI_READ";
        traffic_data[305].size_bytes = 64;
        traffic_data[306].timestamp = 197;
        traffic_data[306].source_node = 6;
        traffic_data[306].dest_node = 14;
        traffic_data[306].packet_type = "CHI_WRITE";
        traffic_data[306].size_bytes = 64;
        traffic_data[307].timestamp = 198;
        traffic_data[307].source_node = 8;
        traffic_data[307].dest_node = 4;
        traffic_data[307].packet_type = "AXI_WRITE";
        traffic_data[307].size_bytes = 64;
        traffic_data[308].timestamp = 200;
        traffic_data[308].source_node = 6;
        traffic_data[308].dest_node = 15;
        traffic_data[308].packet_type = "CHI_READ";
        traffic_data[308].size_bytes = 64;
        traffic_data[309].timestamp = 200;
        traffic_data[309].source_node = 14;
        traffic_data[309].dest_node = 8;
        traffic_data[309].packet_type = "AXI_WRITE";
        traffic_data[309].size_bytes = 64;
        traffic_data[310].timestamp = 201;
        traffic_data[310].source_node = 1;
        traffic_data[310].dest_node = 4;
        traffic_data[310].packet_type = "AXI_WRITE";
        traffic_data[310].size_bytes = 64;
        traffic_data[311].timestamp = 202;
        traffic_data[311].source_node = 1;
        traffic_data[311].dest_node = 15;
        traffic_data[311].packet_type = "CHI_READ";
        traffic_data[311].size_bytes = 64;
        traffic_data[312].timestamp = 202;
        traffic_data[312].source_node = 7;
        traffic_data[312].dest_node = 9;
        traffic_data[312].packet_type = "CHI_READ";
        traffic_data[312].size_bytes = 64;
        traffic_data[313].timestamp = 202;
        traffic_data[313].source_node = 14;
        traffic_data[313].dest_node = 1;
        traffic_data[313].packet_type = "AXI_WRITE";
        traffic_data[313].size_bytes = 64;
        traffic_data[314].timestamp = 203;
        traffic_data[314].source_node = 14;
        traffic_data[314].dest_node = 10;
        traffic_data[314].packet_type = "AXI_WRITE";
        traffic_data[314].size_bytes = 64;
        traffic_data[315].timestamp = 203;
        traffic_data[315].source_node = 15;
        traffic_data[315].dest_node = 11;
        traffic_data[315].packet_type = "CHI_READ";
        traffic_data[315].size_bytes = 64;
        traffic_data[316].timestamp = 204;
        traffic_data[316].source_node = 0;
        traffic_data[316].dest_node = 2;
        traffic_data[316].packet_type = "AXI_READ";
        traffic_data[316].size_bytes = 64;
        traffic_data[317].timestamp = 204;
        traffic_data[317].source_node = 3;
        traffic_data[317].dest_node = 14;
        traffic_data[317].packet_type = "AXI_WRITE";
        traffic_data[317].size_bytes = 64;
        traffic_data[318].timestamp = 204;
        traffic_data[318].source_node = 11;
        traffic_data[318].dest_node = 12;
        traffic_data[318].packet_type = "AXI_READ";
        traffic_data[318].size_bytes = 64;
        traffic_data[319].timestamp = 204;
        traffic_data[319].source_node = 15;
        traffic_data[319].dest_node = 14;
        traffic_data[319].packet_type = "AXI_READ";
        traffic_data[319].size_bytes = 64;
        traffic_data[320].timestamp = 205;
        traffic_data[320].source_node = 7;
        traffic_data[320].dest_node = 2;
        traffic_data[320].packet_type = "AXI_WRITE";
        traffic_data[320].size_bytes = 64;
        traffic_data[321].timestamp = 206;
        traffic_data[321].source_node = 7;
        traffic_data[321].dest_node = 10;
        traffic_data[321].packet_type = "CHI_WRITE";
        traffic_data[321].size_bytes = 64;
        traffic_data[322].timestamp = 207;
        traffic_data[322].source_node = 14;
        traffic_data[322].dest_node = 1;
        traffic_data[322].packet_type = "AXI_WRITE";
        traffic_data[322].size_bytes = 64;
        traffic_data[323].timestamp = 209;
        traffic_data[323].source_node = 0;
        traffic_data[323].dest_node = 4;
        traffic_data[323].packet_type = "AXI_WRITE";
        traffic_data[323].size_bytes = 64;
        traffic_data[324].timestamp = 209;
        traffic_data[324].source_node = 13;
        traffic_data[324].dest_node = 4;
        traffic_data[324].packet_type = "AXI_WRITE";
        traffic_data[324].size_bytes = 64;
        traffic_data[325].timestamp = 210;
        traffic_data[325].source_node = 10;
        traffic_data[325].dest_node = 4;
        traffic_data[325].packet_type = "CHI_WRITE";
        traffic_data[325].size_bytes = 64;
        traffic_data[326].timestamp = 211;
        traffic_data[326].source_node = 3;
        traffic_data[326].dest_node = 6;
        traffic_data[326].packet_type = "AXI_READ";
        traffic_data[326].size_bytes = 64;
        traffic_data[327].timestamp = 212;
        traffic_data[327].source_node = 4;
        traffic_data[327].dest_node = 6;
        traffic_data[327].packet_type = "AXI_WRITE";
        traffic_data[327].size_bytes = 64;
        traffic_data[328].timestamp = 212;
        traffic_data[328].source_node = 5;
        traffic_data[328].dest_node = 3;
        traffic_data[328].packet_type = "CHI_READ";
        traffic_data[328].size_bytes = 64;
        traffic_data[329].timestamp = 212;
        traffic_data[329].source_node = 9;
        traffic_data[329].dest_node = 11;
        traffic_data[329].packet_type = "CHI_READ";
        traffic_data[329].size_bytes = 64;
        traffic_data[330].timestamp = 213;
        traffic_data[330].source_node = 5;
        traffic_data[330].dest_node = 4;
        traffic_data[330].packet_type = "CHI_WRITE";
        traffic_data[330].size_bytes = 64;
        traffic_data[331].timestamp = 213;
        traffic_data[331].source_node = 13;
        traffic_data[331].dest_node = 15;
        traffic_data[331].packet_type = "AXI_WRITE";
        traffic_data[331].size_bytes = 64;
        traffic_data[332].timestamp = 216;
        traffic_data[332].source_node = 15;
        traffic_data[332].dest_node = 6;
        traffic_data[332].packet_type = "CHI_WRITE";
        traffic_data[332].size_bytes = 64;
        traffic_data[333].timestamp = 217;
        traffic_data[333].source_node = 1;
        traffic_data[333].dest_node = 9;
        traffic_data[333].packet_type = "CHI_WRITE";
        traffic_data[333].size_bytes = 64;
        traffic_data[334].timestamp = 217;
        traffic_data[334].source_node = 10;
        traffic_data[334].dest_node = 11;
        traffic_data[334].packet_type = "AXI_WRITE";
        traffic_data[334].size_bytes = 64;
        traffic_data[335].timestamp = 217;
        traffic_data[335].source_node = 13;
        traffic_data[335].dest_node = 12;
        traffic_data[335].packet_type = "CHI_WRITE";
        traffic_data[335].size_bytes = 64;
        traffic_data[336].timestamp = 218;
        traffic_data[336].source_node = 0;
        traffic_data[336].dest_node = 9;
        traffic_data[336].packet_type = "CHI_WRITE";
        traffic_data[336].size_bytes = 64;
        traffic_data[337].timestamp = 218;
        traffic_data[337].source_node = 9;
        traffic_data[337].dest_node = 2;
        traffic_data[337].packet_type = "CHI_READ";
        traffic_data[337].size_bytes = 64;
        traffic_data[338].timestamp = 219;
        traffic_data[338].source_node = 5;
        traffic_data[338].dest_node = 11;
        traffic_data[338].packet_type = "AXI_WRITE";
        traffic_data[338].size_bytes = 64;
        traffic_data[339].timestamp = 221;
        traffic_data[339].source_node = 10;
        traffic_data[339].dest_node = 1;
        traffic_data[339].packet_type = "AXI_WRITE";
        traffic_data[339].size_bytes = 64;
        traffic_data[340].timestamp = 221;
        traffic_data[340].source_node = 13;
        traffic_data[340].dest_node = 4;
        traffic_data[340].packet_type = "AXI_WRITE";
        traffic_data[340].size_bytes = 64;
        traffic_data[341].timestamp = 222;
        traffic_data[341].source_node = 6;
        traffic_data[341].dest_node = 13;
        traffic_data[341].packet_type = "AXI_WRITE";
        traffic_data[341].size_bytes = 64;
        traffic_data[342].timestamp = 222;
        traffic_data[342].source_node = 13;
        traffic_data[342].dest_node = 9;
        traffic_data[342].packet_type = "AXI_WRITE";
        traffic_data[342].size_bytes = 64;
        traffic_data[343].timestamp = 223;
        traffic_data[343].source_node = 3;
        traffic_data[343].dest_node = 5;
        traffic_data[343].packet_type = "CHI_WRITE";
        traffic_data[343].size_bytes = 64;
        traffic_data[344].timestamp = 223;
        traffic_data[344].source_node = 9;
        traffic_data[344].dest_node = 1;
        traffic_data[344].packet_type = "CHI_READ";
        traffic_data[344].size_bytes = 64;
        traffic_data[345].timestamp = 224;
        traffic_data[345].source_node = 3;
        traffic_data[345].dest_node = 2;
        traffic_data[345].packet_type = "CHI_WRITE";
        traffic_data[345].size_bytes = 64;
        traffic_data[346].timestamp = 227;
        traffic_data[346].source_node = 10;
        traffic_data[346].dest_node = 11;
        traffic_data[346].packet_type = "CHI_WRITE";
        traffic_data[346].size_bytes = 64;
        traffic_data[347].timestamp = 227;
        traffic_data[347].source_node = 14;
        traffic_data[347].dest_node = 7;
        traffic_data[347].packet_type = "CHI_READ";
        traffic_data[347].size_bytes = 64;
        traffic_data[348].timestamp = 228;
        traffic_data[348].source_node = 10;
        traffic_data[348].dest_node = 13;
        traffic_data[348].packet_type = "CHI_WRITE";
        traffic_data[348].size_bytes = 64;
        traffic_data[349].timestamp = 229;
        traffic_data[349].source_node = 5;
        traffic_data[349].dest_node = 3;
        traffic_data[349].packet_type = "CHI_WRITE";
        traffic_data[349].size_bytes = 64;
        traffic_data[350].timestamp = 230;
        traffic_data[350].source_node = 9;
        traffic_data[350].dest_node = 4;
        traffic_data[350].packet_type = "AXI_WRITE";
        traffic_data[350].size_bytes = 64;
        traffic_data[351].timestamp = 231;
        traffic_data[351].source_node = 0;
        traffic_data[351].dest_node = 7;
        traffic_data[351].packet_type = "CHI_WRITE";
        traffic_data[351].size_bytes = 64;
        traffic_data[352].timestamp = 231;
        traffic_data[352].source_node = 9;
        traffic_data[352].dest_node = 1;
        traffic_data[352].packet_type = "AXI_WRITE";
        traffic_data[352].size_bytes = 64;
        traffic_data[353].timestamp = 231;
        traffic_data[353].source_node = 10;
        traffic_data[353].dest_node = 14;
        traffic_data[353].packet_type = "CHI_READ";
        traffic_data[353].size_bytes = 64;
        traffic_data[354].timestamp = 232;
        traffic_data[354].source_node = 3;
        traffic_data[354].dest_node = 1;
        traffic_data[354].packet_type = "CHI_READ";
        traffic_data[354].size_bytes = 64;
        traffic_data[355].timestamp = 233;
        traffic_data[355].source_node = 10;
        traffic_data[355].dest_node = 2;
        traffic_data[355].packet_type = "CHI_READ";
        traffic_data[355].size_bytes = 64;
        traffic_data[356].timestamp = 234;
        traffic_data[356].source_node = 8;
        traffic_data[356].dest_node = 12;
        traffic_data[356].packet_type = "AXI_WRITE";
        traffic_data[356].size_bytes = 64;
        traffic_data[357].timestamp = 234;
        traffic_data[357].source_node = 12;
        traffic_data[357].dest_node = 2;
        traffic_data[357].packet_type = "CHI_WRITE";
        traffic_data[357].size_bytes = 64;
        traffic_data[358].timestamp = 234;
        traffic_data[358].source_node = 14;
        traffic_data[358].dest_node = 15;
        traffic_data[358].packet_type = "CHI_WRITE";
        traffic_data[358].size_bytes = 64;
        traffic_data[359].timestamp = 235;
        traffic_data[359].source_node = 0;
        traffic_data[359].dest_node = 7;
        traffic_data[359].packet_type = "AXI_READ";
        traffic_data[359].size_bytes = 64;
        traffic_data[360].timestamp = 235;
        traffic_data[360].source_node = 3;
        traffic_data[360].dest_node = 15;
        traffic_data[360].packet_type = "CHI_WRITE";
        traffic_data[360].size_bytes = 64;
        traffic_data[361].timestamp = 235;
        traffic_data[361].source_node = 10;
        traffic_data[361].dest_node = 11;
        traffic_data[361].packet_type = "CHI_READ";
        traffic_data[361].size_bytes = 64;
        traffic_data[362].timestamp = 237;
        traffic_data[362].source_node = 3;
        traffic_data[362].dest_node = 14;
        traffic_data[362].packet_type = "AXI_WRITE";
        traffic_data[362].size_bytes = 64;
        traffic_data[363].timestamp = 237;
        traffic_data[363].source_node = 6;
        traffic_data[363].dest_node = 15;
        traffic_data[363].packet_type = "CHI_WRITE";
        traffic_data[363].size_bytes = 64;
        traffic_data[364].timestamp = 237;
        traffic_data[364].source_node = 9;
        traffic_data[364].dest_node = 6;
        traffic_data[364].packet_type = "CHI_READ";
        traffic_data[364].size_bytes = 64;
        traffic_data[365].timestamp = 238;
        traffic_data[365].source_node = 5;
        traffic_data[365].dest_node = 11;
        traffic_data[365].packet_type = "AXI_WRITE";
        traffic_data[365].size_bytes = 64;
        traffic_data[366].timestamp = 238;
        traffic_data[366].source_node = 15;
        traffic_data[366].dest_node = 2;
        traffic_data[366].packet_type = "CHI_READ";
        traffic_data[366].size_bytes = 64;
        traffic_data[367].timestamp = 239;
        traffic_data[367].source_node = 8;
        traffic_data[367].dest_node = 1;
        traffic_data[367].packet_type = "CHI_READ";
        traffic_data[367].size_bytes = 64;
        traffic_data[368].timestamp = 240;
        traffic_data[368].source_node = 8;
        traffic_data[368].dest_node = 13;
        traffic_data[368].packet_type = "CHI_WRITE";
        traffic_data[368].size_bytes = 64;
        traffic_data[369].timestamp = 240;
        traffic_data[369].source_node = 9;
        traffic_data[369].dest_node = 7;
        traffic_data[369].packet_type = "AXI_WRITE";
        traffic_data[369].size_bytes = 64;
        traffic_data[370].timestamp = 241;
        traffic_data[370].source_node = 4;
        traffic_data[370].dest_node = 8;
        traffic_data[370].packet_type = "AXI_READ";
        traffic_data[370].size_bytes = 64;
        traffic_data[371].timestamp = 241;
        traffic_data[371].source_node = 12;
        traffic_data[371].dest_node = 15;
        traffic_data[371].packet_type = "AXI_READ";
        traffic_data[371].size_bytes = 64;
        traffic_data[372].timestamp = 242;
        traffic_data[372].source_node = 10;
        traffic_data[372].dest_node = 0;
        traffic_data[372].packet_type = "CHI_WRITE";
        traffic_data[372].size_bytes = 64;
        traffic_data[373].timestamp = 243;
        traffic_data[373].source_node = 4;
        traffic_data[373].dest_node = 6;
        traffic_data[373].packet_type = "AXI_WRITE";
        traffic_data[373].size_bytes = 64;
        traffic_data[374].timestamp = 244;
        traffic_data[374].source_node = 15;
        traffic_data[374].dest_node = 2;
        traffic_data[374].packet_type = "CHI_WRITE";
        traffic_data[374].size_bytes = 64;
        traffic_data[375].timestamp = 245;
        traffic_data[375].source_node = 3;
        traffic_data[375].dest_node = 11;
        traffic_data[375].packet_type = "CHI_WRITE";
        traffic_data[375].size_bytes = 64;
        traffic_data[376].timestamp = 245;
        traffic_data[376].source_node = 10;
        traffic_data[376].dest_node = 8;
        traffic_data[376].packet_type = "CHI_WRITE";
        traffic_data[376].size_bytes = 64;
        traffic_data[377].timestamp = 246;
        traffic_data[377].source_node = 2;
        traffic_data[377].dest_node = 11;
        traffic_data[377].packet_type = "AXI_READ";
        traffic_data[377].size_bytes = 64;
        traffic_data[378].timestamp = 246;
        traffic_data[378].source_node = 3;
        traffic_data[378].dest_node = 2;
        traffic_data[378].packet_type = "AXI_WRITE";
        traffic_data[378].size_bytes = 64;
        traffic_data[379].timestamp = 246;
        traffic_data[379].source_node = 7;
        traffic_data[379].dest_node = 10;
        traffic_data[379].packet_type = "CHI_WRITE";
        traffic_data[379].size_bytes = 64;
        traffic_data[380].timestamp = 246;
        traffic_data[380].source_node = 14;
        traffic_data[380].dest_node = 15;
        traffic_data[380].packet_type = "AXI_WRITE";
        traffic_data[380].size_bytes = 64;
        traffic_data[381].timestamp = 247;
        traffic_data[381].source_node = 9;
        traffic_data[381].dest_node = 10;
        traffic_data[381].packet_type = "CHI_READ";
        traffic_data[381].size_bytes = 64;
        traffic_data[382].timestamp = 247;
        traffic_data[382].source_node = 13;
        traffic_data[382].dest_node = 3;
        traffic_data[382].packet_type = "AXI_READ";
        traffic_data[382].size_bytes = 64;
        traffic_data[383].timestamp = 250;
        traffic_data[383].source_node = 5;
        traffic_data[383].dest_node = 0;
        traffic_data[383].packet_type = "CHI_READ";
        traffic_data[383].size_bytes = 64;
        traffic_data[384].timestamp = 250;
        traffic_data[384].source_node = 13;
        traffic_data[384].dest_node = 14;
        traffic_data[384].packet_type = "CHI_READ";
        traffic_data[384].size_bytes = 64;
        traffic_data[385].timestamp = 251;
        traffic_data[385].source_node = 2;
        traffic_data[385].dest_node = 8;
        traffic_data[385].packet_type = "CHI_READ";
        traffic_data[385].size_bytes = 64;
        traffic_data[386].timestamp = 251;
        traffic_data[386].source_node = 12;
        traffic_data[386].dest_node = 5;
        traffic_data[386].packet_type = "CHI_WRITE";
        traffic_data[386].size_bytes = 64;
        traffic_data[387].timestamp = 252;
        traffic_data[387].source_node = 6;
        traffic_data[387].dest_node = 0;
        traffic_data[387].packet_type = "CHI_READ";
        traffic_data[387].size_bytes = 64;
        traffic_data[388].timestamp = 252;
        traffic_data[388].source_node = 15;
        traffic_data[388].dest_node = 12;
        traffic_data[388].packet_type = "CHI_WRITE";
        traffic_data[388].size_bytes = 64;
        traffic_data[389].timestamp = 253;
        traffic_data[389].source_node = 0;
        traffic_data[389].dest_node = 9;
        traffic_data[389].packet_type = "AXI_READ";
        traffic_data[389].size_bytes = 64;
        traffic_data[390].timestamp = 253;
        traffic_data[390].source_node = 11;
        traffic_data[390].dest_node = 6;
        traffic_data[390].packet_type = "CHI_READ";
        traffic_data[390].size_bytes = 64;
        traffic_data[391].timestamp = 256;
        traffic_data[391].source_node = 5;
        traffic_data[391].dest_node = 12;
        traffic_data[391].packet_type = "AXI_READ";
        traffic_data[391].size_bytes = 64;
        traffic_data[392].timestamp = 257;
        traffic_data[392].source_node = 13;
        traffic_data[392].dest_node = 3;
        traffic_data[392].packet_type = "CHI_READ";
        traffic_data[392].size_bytes = 64;
        traffic_data[393].timestamp = 257;
        traffic_data[393].source_node = 14;
        traffic_data[393].dest_node = 10;
        traffic_data[393].packet_type = "AXI_READ";
        traffic_data[393].size_bytes = 64;
        traffic_data[394].timestamp = 257;
        traffic_data[394].source_node = 15;
        traffic_data[394].dest_node = 10;
        traffic_data[394].packet_type = "CHI_READ";
        traffic_data[394].size_bytes = 64;
        traffic_data[395].timestamp = 258;
        traffic_data[395].source_node = 13;
        traffic_data[395].dest_node = 3;
        traffic_data[395].packet_type = "CHI_WRITE";
        traffic_data[395].size_bytes = 64;
        traffic_data[396].timestamp = 259;
        traffic_data[396].source_node = 0;
        traffic_data[396].dest_node = 15;
        traffic_data[396].packet_type = "CHI_READ";
        traffic_data[396].size_bytes = 64;
        traffic_data[397].timestamp = 259;
        traffic_data[397].source_node = 15;
        traffic_data[397].dest_node = 8;
        traffic_data[397].packet_type = "CHI_READ";
        traffic_data[397].size_bytes = 64;
        traffic_data[398].timestamp = 261;
        traffic_data[398].source_node = 14;
        traffic_data[398].dest_node = 8;
        traffic_data[398].packet_type = "AXI_READ";
        traffic_data[398].size_bytes = 64;
        traffic_data[399].timestamp = 262;
        traffic_data[399].source_node = 2;
        traffic_data[399].dest_node = 6;
        traffic_data[399].packet_type = "CHI_WRITE";
        traffic_data[399].size_bytes = 64;
        traffic_data[400].timestamp = 262;
        traffic_data[400].source_node = 12;
        traffic_data[400].dest_node = 9;
        traffic_data[400].packet_type = "CHI_READ";
        traffic_data[400].size_bytes = 64;
        traffic_data[401].timestamp = 263;
        traffic_data[401].source_node = 1;
        traffic_data[401].dest_node = 2;
        traffic_data[401].packet_type = "CHI_WRITE";
        traffic_data[401].size_bytes = 64;
        traffic_data[402].timestamp = 265;
        traffic_data[402].source_node = 5;
        traffic_data[402].dest_node = 1;
        traffic_data[402].packet_type = "CHI_WRITE";
        traffic_data[402].size_bytes = 64;
        traffic_data[403].timestamp = 265;
        traffic_data[403].source_node = 12;
        traffic_data[403].dest_node = 6;
        traffic_data[403].packet_type = "AXI_READ";
        traffic_data[403].size_bytes = 64;
        traffic_data[404].timestamp = 266;
        traffic_data[404].source_node = 9;
        traffic_data[404].dest_node = 8;
        traffic_data[404].packet_type = "AXI_READ";
        traffic_data[404].size_bytes = 64;
        traffic_data[405].timestamp = 267;
        traffic_data[405].source_node = 0;
        traffic_data[405].dest_node = 8;
        traffic_data[405].packet_type = "AXI_WRITE";
        traffic_data[405].size_bytes = 64;
        traffic_data[406].timestamp = 267;
        traffic_data[406].source_node = 2;
        traffic_data[406].dest_node = 6;
        traffic_data[406].packet_type = "AXI_WRITE";
        traffic_data[406].size_bytes = 64;
        traffic_data[407].timestamp = 269;
        traffic_data[407].source_node = 4;
        traffic_data[407].dest_node = 15;
        traffic_data[407].packet_type = "CHI_WRITE";
        traffic_data[407].size_bytes = 64;
        traffic_data[408].timestamp = 269;
        traffic_data[408].source_node = 9;
        traffic_data[408].dest_node = 10;
        traffic_data[408].packet_type = "AXI_READ";
        traffic_data[408].size_bytes = 64;
        traffic_data[409].timestamp = 269;
        traffic_data[409].source_node = 15;
        traffic_data[409].dest_node = 2;
        traffic_data[409].packet_type = "AXI_READ";
        traffic_data[409].size_bytes = 64;
        traffic_data[410].timestamp = 270;
        traffic_data[410].source_node = 1;
        traffic_data[410].dest_node = 14;
        traffic_data[410].packet_type = "AXI_READ";
        traffic_data[410].size_bytes = 64;
        traffic_data[411].timestamp = 270;
        traffic_data[411].source_node = 6;
        traffic_data[411].dest_node = 7;
        traffic_data[411].packet_type = "AXI_WRITE";
        traffic_data[411].size_bytes = 64;
        traffic_data[412].timestamp = 271;
        traffic_data[412].source_node = 0;
        traffic_data[412].dest_node = 13;
        traffic_data[412].packet_type = "CHI_READ";
        traffic_data[412].size_bytes = 64;
        traffic_data[413].timestamp = 271;
        traffic_data[413].source_node = 6;
        traffic_data[413].dest_node = 8;
        traffic_data[413].packet_type = "AXI_WRITE";
        traffic_data[413].size_bytes = 64;
        traffic_data[414].timestamp = 271;
        traffic_data[414].source_node = 13;
        traffic_data[414].dest_node = 9;
        traffic_data[414].packet_type = "AXI_READ";
        traffic_data[414].size_bytes = 64;
        traffic_data[415].timestamp = 273;
        traffic_data[415].source_node = 1;
        traffic_data[415].dest_node = 0;
        traffic_data[415].packet_type = "CHI_WRITE";
        traffic_data[415].size_bytes = 64;
        traffic_data[416].timestamp = 273;
        traffic_data[416].source_node = 11;
        traffic_data[416].dest_node = 3;
        traffic_data[416].packet_type = "CHI_READ";
        traffic_data[416].size_bytes = 64;
        traffic_data[417].timestamp = 273;
        traffic_data[417].source_node = 13;
        traffic_data[417].dest_node = 4;
        traffic_data[417].packet_type = "CHI_READ";
        traffic_data[417].size_bytes = 64;
        traffic_data[418].timestamp = 274;
        traffic_data[418].source_node = 10;
        traffic_data[418].dest_node = 2;
        traffic_data[418].packet_type = "CHI_WRITE";
        traffic_data[418].size_bytes = 64;
        traffic_data[419].timestamp = 275;
        traffic_data[419].source_node = 2;
        traffic_data[419].dest_node = 9;
        traffic_data[419].packet_type = "CHI_READ";
        traffic_data[419].size_bytes = 64;
        traffic_data[420].timestamp = 275;
        traffic_data[420].source_node = 6;
        traffic_data[420].dest_node = 10;
        traffic_data[420].packet_type = "CHI_READ";
        traffic_data[420].size_bytes = 64;
        traffic_data[421].timestamp = 275;
        traffic_data[421].source_node = 12;
        traffic_data[421].dest_node = 6;
        traffic_data[421].packet_type = "AXI_WRITE";
        traffic_data[421].size_bytes = 64;
        traffic_data[422].timestamp = 276;
        traffic_data[422].source_node = 4;
        traffic_data[422].dest_node = 7;
        traffic_data[422].packet_type = "AXI_READ";
        traffic_data[422].size_bytes = 64;
        traffic_data[423].timestamp = 277;
        traffic_data[423].source_node = 0;
        traffic_data[423].dest_node = 8;
        traffic_data[423].packet_type = "AXI_WRITE";
        traffic_data[423].size_bytes = 64;
        traffic_data[424].timestamp = 278;
        traffic_data[424].source_node = 0;
        traffic_data[424].dest_node = 15;
        traffic_data[424].packet_type = "AXI_READ";
        traffic_data[424].size_bytes = 64;
        traffic_data[425].timestamp = 278;
        traffic_data[425].source_node = 3;
        traffic_data[425].dest_node = 8;
        traffic_data[425].packet_type = "AXI_READ";
        traffic_data[425].size_bytes = 64;
        traffic_data[426].timestamp = 278;
        traffic_data[426].source_node = 7;
        traffic_data[426].dest_node = 13;
        traffic_data[426].packet_type = "CHI_READ";
        traffic_data[426].size_bytes = 64;
        traffic_data[427].timestamp = 279;
        traffic_data[427].source_node = 15;
        traffic_data[427].dest_node = 0;
        traffic_data[427].packet_type = "CHI_WRITE";
        traffic_data[427].size_bytes = 64;
        traffic_data[428].timestamp = 280;
        traffic_data[428].source_node = 1;
        traffic_data[428].dest_node = 7;
        traffic_data[428].packet_type = "AXI_READ";
        traffic_data[428].size_bytes = 64;
        traffic_data[429].timestamp = 280;
        traffic_data[429].source_node = 2;
        traffic_data[429].dest_node = 7;
        traffic_data[429].packet_type = "AXI_WRITE";
        traffic_data[429].size_bytes = 64;
        traffic_data[430].timestamp = 280;
        traffic_data[430].source_node = 13;
        traffic_data[430].dest_node = 15;
        traffic_data[430].packet_type = "CHI_WRITE";
        traffic_data[430].size_bytes = 64;
        traffic_data[431].timestamp = 280;
        traffic_data[431].source_node = 15;
        traffic_data[431].dest_node = 12;
        traffic_data[431].packet_type = "CHI_WRITE";
        traffic_data[431].size_bytes = 64;
        traffic_data[432].timestamp = 281;
        traffic_data[432].source_node = 0;
        traffic_data[432].dest_node = 5;
        traffic_data[432].packet_type = "CHI_WRITE";
        traffic_data[432].size_bytes = 64;
        traffic_data[433].timestamp = 281;
        traffic_data[433].source_node = 13;
        traffic_data[433].dest_node = 1;
        traffic_data[433].packet_type = "CHI_READ";
        traffic_data[433].size_bytes = 64;
        traffic_data[434].timestamp = 282;
        traffic_data[434].source_node = 8;
        traffic_data[434].dest_node = 4;
        traffic_data[434].packet_type = "CHI_WRITE";
        traffic_data[434].size_bytes = 64;
        traffic_data[435].timestamp = 283;
        traffic_data[435].source_node = 8;
        traffic_data[435].dest_node = 15;
        traffic_data[435].packet_type = "CHI_WRITE";
        traffic_data[435].size_bytes = 64;
        traffic_data[436].timestamp = 283;
        traffic_data[436].source_node = 12;
        traffic_data[436].dest_node = 7;
        traffic_data[436].packet_type = "AXI_WRITE";
        traffic_data[436].size_bytes = 64;
        traffic_data[437].timestamp = 284;
        traffic_data[437].source_node = 5;
        traffic_data[437].dest_node = 3;
        traffic_data[437].packet_type = "AXI_WRITE";
        traffic_data[437].size_bytes = 64;
        traffic_data[438].timestamp = 284;
        traffic_data[438].source_node = 9;
        traffic_data[438].dest_node = 2;
        traffic_data[438].packet_type = "AXI_WRITE";
        traffic_data[438].size_bytes = 64;
        traffic_data[439].timestamp = 285;
        traffic_data[439].source_node = 13;
        traffic_data[439].dest_node = 15;
        traffic_data[439].packet_type = "AXI_READ";
        traffic_data[439].size_bytes = 64;
        traffic_data[440].timestamp = 285;
        traffic_data[440].source_node = 14;
        traffic_data[440].dest_node = 8;
        traffic_data[440].packet_type = "CHI_READ";
        traffic_data[440].size_bytes = 64;
        traffic_data[441].timestamp = 286;
        traffic_data[441].source_node = 1;
        traffic_data[441].dest_node = 7;
        traffic_data[441].packet_type = "CHI_WRITE";
        traffic_data[441].size_bytes = 64;
        traffic_data[442].timestamp = 287;
        traffic_data[442].source_node = 0;
        traffic_data[442].dest_node = 11;
        traffic_data[442].packet_type = "AXI_READ";
        traffic_data[442].size_bytes = 64;
        traffic_data[443].timestamp = 288;
        traffic_data[443].source_node = 3;
        traffic_data[443].dest_node = 8;
        traffic_data[443].packet_type = "AXI_WRITE";
        traffic_data[443].size_bytes = 64;
        traffic_data[444].timestamp = 288;
        traffic_data[444].source_node = 8;
        traffic_data[444].dest_node = 0;
        traffic_data[444].packet_type = "CHI_WRITE";
        traffic_data[444].size_bytes = 64;
        traffic_data[445].timestamp = 289;
        traffic_data[445].source_node = 3;
        traffic_data[445].dest_node = 15;
        traffic_data[445].packet_type = "AXI_READ";
        traffic_data[445].size_bytes = 64;
        traffic_data[446].timestamp = 289;
        traffic_data[446].source_node = 14;
        traffic_data[446].dest_node = 7;
        traffic_data[446].packet_type = "CHI_WRITE";
        traffic_data[446].size_bytes = 64;
        traffic_data[447].timestamp = 291;
        traffic_data[447].source_node = 0;
        traffic_data[447].dest_node = 8;
        traffic_data[447].packet_type = "AXI_READ";
        traffic_data[447].size_bytes = 64;
        traffic_data[448].timestamp = 291;
        traffic_data[448].source_node = 2;
        traffic_data[448].dest_node = 13;
        traffic_data[448].packet_type = "CHI_READ";
        traffic_data[448].size_bytes = 64;
        traffic_data[449].timestamp = 292;
        traffic_data[449].source_node = 2;
        traffic_data[449].dest_node = 1;
        traffic_data[449].packet_type = "AXI_WRITE";
        traffic_data[449].size_bytes = 64;
        traffic_data[450].timestamp = 292;
        traffic_data[450].source_node = 14;
        traffic_data[450].dest_node = 4;
        traffic_data[450].packet_type = "AXI_READ";
        traffic_data[450].size_bytes = 64;
        traffic_data[451].timestamp = 292;
        traffic_data[451].source_node = 15;
        traffic_data[451].dest_node = 7;
        traffic_data[451].packet_type = "CHI_WRITE";
        traffic_data[451].size_bytes = 64;
        traffic_data[452].timestamp = 294;
        traffic_data[452].source_node = 0;
        traffic_data[452].dest_node = 9;
        traffic_data[452].packet_type = "CHI_READ";
        traffic_data[452].size_bytes = 64;
        traffic_data[453].timestamp = 294;
        traffic_data[453].source_node = 7;
        traffic_data[453].dest_node = 11;
        traffic_data[453].packet_type = "CHI_WRITE";
        traffic_data[453].size_bytes = 64;
        traffic_data[454].timestamp = 295;
        traffic_data[454].source_node = 1;
        traffic_data[454].dest_node = 0;
        traffic_data[454].packet_type = "AXI_READ";
        traffic_data[454].size_bytes = 64;
        traffic_data[455].timestamp = 295;
        traffic_data[455].source_node = 2;
        traffic_data[455].dest_node = 1;
        traffic_data[455].packet_type = "AXI_READ";
        traffic_data[455].size_bytes = 64;
        traffic_data[456].timestamp = 295;
        traffic_data[456].source_node = 7;
        traffic_data[456].dest_node = 10;
        traffic_data[456].packet_type = "AXI_READ";
        traffic_data[456].size_bytes = 64;
        traffic_data[457].timestamp = 295;
        traffic_data[457].source_node = 8;
        traffic_data[457].dest_node = 10;
        traffic_data[457].packet_type = "AXI_WRITE";
        traffic_data[457].size_bytes = 64;
        traffic_data[458].timestamp = 297;
        traffic_data[458].source_node = 0;
        traffic_data[458].dest_node = 13;
        traffic_data[458].packet_type = "AXI_READ";
        traffic_data[458].size_bytes = 64;
        traffic_data[459].timestamp = 297;
        traffic_data[459].source_node = 3;
        traffic_data[459].dest_node = 14;
        traffic_data[459].packet_type = "CHI_READ";
        traffic_data[459].size_bytes = 64;
        traffic_data[460].timestamp = 297;
        traffic_data[460].source_node = 5;
        traffic_data[460].dest_node = 15;
        traffic_data[460].packet_type = "AXI_WRITE";
        traffic_data[460].size_bytes = 64;
        traffic_data[461].timestamp = 298;
        traffic_data[461].source_node = 0;
        traffic_data[461].dest_node = 10;
        traffic_data[461].packet_type = "CHI_READ";
        traffic_data[461].size_bytes = 64;
        traffic_data[462].timestamp = 298;
        traffic_data[462].source_node = 2;
        traffic_data[462].dest_node = 8;
        traffic_data[462].packet_type = "AXI_WRITE";
        traffic_data[462].size_bytes = 64;
        traffic_data[463].timestamp = 298;
        traffic_data[463].source_node = 4;
        traffic_data[463].dest_node = 0;
        traffic_data[463].packet_type = "CHI_WRITE";
        traffic_data[463].size_bytes = 64;
        traffic_data[464].timestamp = 299;
        traffic_data[464].source_node = 1;
        traffic_data[464].dest_node = 12;
        traffic_data[464].packet_type = "CHI_WRITE";
        traffic_data[464].size_bytes = 64;
        traffic_data[465].timestamp = 299;
        traffic_data[465].source_node = 7;
        traffic_data[465].dest_node = 11;
        traffic_data[465].packet_type = "AXI_READ";
        traffic_data[465].size_bytes = 64;
        traffic_data[466].timestamp = 300;
        traffic_data[466].source_node = 10;
        traffic_data[466].dest_node = 0;
        traffic_data[466].packet_type = "AXI_WRITE";
        traffic_data[466].size_bytes = 64;
        traffic_data[467].timestamp = 300;
        traffic_data[467].source_node = 12;
        traffic_data[467].dest_node = 8;
        traffic_data[467].packet_type = "CHI_READ";
        traffic_data[467].size_bytes = 64;
        traffic_data[468].timestamp = 301;
        traffic_data[468].source_node = 1;
        traffic_data[468].dest_node = 6;
        traffic_data[468].packet_type = "AXI_READ";
        traffic_data[468].size_bytes = 64;
        traffic_data[469].timestamp = 301;
        traffic_data[469].source_node = 13;
        traffic_data[469].dest_node = 11;
        traffic_data[469].packet_type = "AXI_WRITE";
        traffic_data[469].size_bytes = 64;
        traffic_data[470].timestamp = 301;
        traffic_data[470].source_node = 15;
        traffic_data[470].dest_node = 14;
        traffic_data[470].packet_type = "AXI_READ";
        traffic_data[470].size_bytes = 64;
        traffic_data[471].timestamp = 302;
        traffic_data[471].source_node = 2;
        traffic_data[471].dest_node = 11;
        traffic_data[471].packet_type = "AXI_READ";
        traffic_data[471].size_bytes = 64;
        traffic_data[472].timestamp = 302;
        traffic_data[472].source_node = 5;
        traffic_data[472].dest_node = 10;
        traffic_data[472].packet_type = "AXI_WRITE";
        traffic_data[472].size_bytes = 64;
        traffic_data[473].timestamp = 302;
        traffic_data[473].source_node = 7;
        traffic_data[473].dest_node = 14;
        traffic_data[473].packet_type = "AXI_READ";
        traffic_data[473].size_bytes = 64;
        traffic_data[474].timestamp = 302;
        traffic_data[474].source_node = 11;
        traffic_data[474].dest_node = 3;
        traffic_data[474].packet_type = "CHI_WRITE";
        traffic_data[474].size_bytes = 64;
        traffic_data[475].timestamp = 303;
        traffic_data[475].source_node = 6;
        traffic_data[475].dest_node = 2;
        traffic_data[475].packet_type = "CHI_READ";
        traffic_data[475].size_bytes = 64;
        traffic_data[476].timestamp = 303;
        traffic_data[476].source_node = 7;
        traffic_data[476].dest_node = 4;
        traffic_data[476].packet_type = "AXI_WRITE";
        traffic_data[476].size_bytes = 64;
        traffic_data[477].timestamp = 304;
        traffic_data[477].source_node = 4;
        traffic_data[477].dest_node = 0;
        traffic_data[477].packet_type = "AXI_WRITE";
        traffic_data[477].size_bytes = 64;
        traffic_data[478].timestamp = 305;
        traffic_data[478].source_node = 6;
        traffic_data[478].dest_node = 14;
        traffic_data[478].packet_type = "CHI_READ";
        traffic_data[478].size_bytes = 64;
        traffic_data[479].timestamp = 305;
        traffic_data[479].source_node = 8;
        traffic_data[479].dest_node = 3;
        traffic_data[479].packet_type = "AXI_WRITE";
        traffic_data[479].size_bytes = 64;
        traffic_data[480].timestamp = 305;
        traffic_data[480].source_node = 11;
        traffic_data[480].dest_node = 5;
        traffic_data[480].packet_type = "AXI_WRITE";
        traffic_data[480].size_bytes = 64;
        traffic_data[481].timestamp = 305;
        traffic_data[481].source_node = 15;
        traffic_data[481].dest_node = 1;
        traffic_data[481].packet_type = "AXI_WRITE";
        traffic_data[481].size_bytes = 64;
        traffic_data[482].timestamp = 306;
        traffic_data[482].source_node = 5;
        traffic_data[482].dest_node = 11;
        traffic_data[482].packet_type = "CHI_READ";
        traffic_data[482].size_bytes = 64;
        traffic_data[483].timestamp = 306;
        traffic_data[483].source_node = 11;
        traffic_data[483].dest_node = 12;
        traffic_data[483].packet_type = "AXI_READ";
        traffic_data[483].size_bytes = 64;
        traffic_data[484].timestamp = 307;
        traffic_data[484].source_node = 10;
        traffic_data[484].dest_node = 12;
        traffic_data[484].packet_type = "CHI_WRITE";
        traffic_data[484].size_bytes = 64;
        traffic_data[485].timestamp = 308;
        traffic_data[485].source_node = 12;
        traffic_data[485].dest_node = 2;
        traffic_data[485].packet_type = "AXI_READ";
        traffic_data[485].size_bytes = 64;
        traffic_data[486].timestamp = 309;
        traffic_data[486].source_node = 9;
        traffic_data[486].dest_node = 14;
        traffic_data[486].packet_type = "CHI_WRITE";
        traffic_data[486].size_bytes = 64;
        traffic_data[487].timestamp = 309;
        traffic_data[487].source_node = 14;
        traffic_data[487].dest_node = 6;
        traffic_data[487].packet_type = "AXI_WRITE";
        traffic_data[487].size_bytes = 64;
        traffic_data[488].timestamp = 310;
        traffic_data[488].source_node = 7;
        traffic_data[488].dest_node = 8;
        traffic_data[488].packet_type = "AXI_READ";
        traffic_data[488].size_bytes = 64;
        traffic_data[489].timestamp = 310;
        traffic_data[489].source_node = 12;
        traffic_data[489].dest_node = 7;
        traffic_data[489].packet_type = "AXI_WRITE";
        traffic_data[489].size_bytes = 64;
        traffic_data[490].timestamp = 310;
        traffic_data[490].source_node = 13;
        traffic_data[490].dest_node = 12;
        traffic_data[490].packet_type = "AXI_READ";
        traffic_data[490].size_bytes = 64;
        traffic_data[491].timestamp = 311;
        traffic_data[491].source_node = 4;
        traffic_data[491].dest_node = 11;
        traffic_data[491].packet_type = "CHI_READ";
        traffic_data[491].size_bytes = 64;
        traffic_data[492].timestamp = 312;
        traffic_data[492].source_node = 1;
        traffic_data[492].dest_node = 11;
        traffic_data[492].packet_type = "AXI_READ";
        traffic_data[492].size_bytes = 64;
        traffic_data[493].timestamp = 313;
        traffic_data[493].source_node = 2;
        traffic_data[493].dest_node = 7;
        traffic_data[493].packet_type = "CHI_READ";
        traffic_data[493].size_bytes = 64;
        traffic_data[494].timestamp = 313;
        traffic_data[494].source_node = 4;
        traffic_data[494].dest_node = 6;
        traffic_data[494].packet_type = "AXI_WRITE";
        traffic_data[494].size_bytes = 64;
        traffic_data[495].timestamp = 314;
        traffic_data[495].source_node = 7;
        traffic_data[495].dest_node = 5;
        traffic_data[495].packet_type = "CHI_READ";
        traffic_data[495].size_bytes = 64;
        traffic_data[496].timestamp = 315;
        traffic_data[496].source_node = 7;
        traffic_data[496].dest_node = 6;
        traffic_data[496].packet_type = "AXI_WRITE";
        traffic_data[496].size_bytes = 64;
        traffic_data[497].timestamp = 316;
        traffic_data[497].source_node = 9;
        traffic_data[497].dest_node = 14;
        traffic_data[497].packet_type = "AXI_WRITE";
        traffic_data[497].size_bytes = 64;
        traffic_data[498].timestamp = 319;
        traffic_data[498].source_node = 7;
        traffic_data[498].dest_node = 15;
        traffic_data[498].packet_type = "CHI_WRITE";
        traffic_data[498].size_bytes = 64;
        traffic_data[499].timestamp = 320;
        traffic_data[499].source_node = 12;
        traffic_data[499].dest_node = 10;
        traffic_data[499].packet_type = "AXI_READ";
        traffic_data[499].size_bytes = 64;
        traffic_data[500].timestamp = 321;
        traffic_data[500].source_node = 1;
        traffic_data[500].dest_node = 0;
        traffic_data[500].packet_type = "AXI_WRITE";
        traffic_data[500].size_bytes = 64;
        traffic_data[501].timestamp = 321;
        traffic_data[501].source_node = 6;
        traffic_data[501].dest_node = 9;
        traffic_data[501].packet_type = "CHI_WRITE";
        traffic_data[501].size_bytes = 64;
        traffic_data[502].timestamp = 321;
        traffic_data[502].source_node = 14;
        traffic_data[502].dest_node = 10;
        traffic_data[502].packet_type = "CHI_READ";
        traffic_data[502].size_bytes = 64;
        traffic_data[503].timestamp = 322;
        traffic_data[503].source_node = 3;
        traffic_data[503].dest_node = 6;
        traffic_data[503].packet_type = "CHI_READ";
        traffic_data[503].size_bytes = 64;
        traffic_data[504].timestamp = 323;
        traffic_data[504].source_node = 11;
        traffic_data[504].dest_node = 10;
        traffic_data[504].packet_type = "CHI_READ";
        traffic_data[504].size_bytes = 64;
        traffic_data[505].timestamp = 324;
        traffic_data[505].source_node = 4;
        traffic_data[505].dest_node = 14;
        traffic_data[505].packet_type = "CHI_READ";
        traffic_data[505].size_bytes = 64;
        traffic_data[506].timestamp = 324;
        traffic_data[506].source_node = 9;
        traffic_data[506].dest_node = 0;
        traffic_data[506].packet_type = "AXI_WRITE";
        traffic_data[506].size_bytes = 64;
        traffic_data[507].timestamp = 325;
        traffic_data[507].source_node = 7;
        traffic_data[507].dest_node = 12;
        traffic_data[507].packet_type = "CHI_READ";
        traffic_data[507].size_bytes = 64;
        traffic_data[508].timestamp = 326;
        traffic_data[508].source_node = 3;
        traffic_data[508].dest_node = 6;
        traffic_data[508].packet_type = "CHI_WRITE";
        traffic_data[508].size_bytes = 64;
        traffic_data[509].timestamp = 327;
        traffic_data[509].source_node = 1;
        traffic_data[509].dest_node = 13;
        traffic_data[509].packet_type = "AXI_WRITE";
        traffic_data[509].size_bytes = 64;
        traffic_data[510].timestamp = 327;
        traffic_data[510].source_node = 9;
        traffic_data[510].dest_node = 10;
        traffic_data[510].packet_type = "CHI_READ";
        traffic_data[510].size_bytes = 64;
        traffic_data[511].timestamp = 327;
        traffic_data[511].source_node = 11;
        traffic_data[511].dest_node = 8;
        traffic_data[511].packet_type = "CHI_READ";
        traffic_data[511].size_bytes = 64;
        traffic_data[512].timestamp = 328;
        traffic_data[512].source_node = 13;
        traffic_data[512].dest_node = 14;
        traffic_data[512].packet_type = "AXI_WRITE";
        traffic_data[512].size_bytes = 64;
        traffic_data[513].timestamp = 329;
        traffic_data[513].source_node = 8;
        traffic_data[513].dest_node = 14;
        traffic_data[513].packet_type = "AXI_READ";
        traffic_data[513].size_bytes = 64;
        traffic_data[514].timestamp = 329;
        traffic_data[514].source_node = 15;
        traffic_data[514].dest_node = 11;
        traffic_data[514].packet_type = "AXI_READ";
        traffic_data[514].size_bytes = 64;
        traffic_data[515].timestamp = 330;
        traffic_data[515].source_node = 0;
        traffic_data[515].dest_node = 13;
        traffic_data[515].packet_type = "CHI_WRITE";
        traffic_data[515].size_bytes = 64;
        traffic_data[516].timestamp = 330;
        traffic_data[516].source_node = 2;
        traffic_data[516].dest_node = 1;
        traffic_data[516].packet_type = "AXI_READ";
        traffic_data[516].size_bytes = 64;
        traffic_data[517].timestamp = 330;
        traffic_data[517].source_node = 5;
        traffic_data[517].dest_node = 1;
        traffic_data[517].packet_type = "CHI_READ";
        traffic_data[517].size_bytes = 64;
        traffic_data[518].timestamp = 330;
        traffic_data[518].source_node = 6;
        traffic_data[518].dest_node = 4;
        traffic_data[518].packet_type = "AXI_READ";
        traffic_data[518].size_bytes = 64;
        traffic_data[519].timestamp = 330;
        traffic_data[519].source_node = 14;
        traffic_data[519].dest_node = 13;
        traffic_data[519].packet_type = "CHI_READ";
        traffic_data[519].size_bytes = 64;
        traffic_data[520].timestamp = 331;
        traffic_data[520].source_node = 6;
        traffic_data[520].dest_node = 10;
        traffic_data[520].packet_type = "AXI_READ";
        traffic_data[520].size_bytes = 64;
        traffic_data[521].timestamp = 331;
        traffic_data[521].source_node = 12;
        traffic_data[521].dest_node = 11;
        traffic_data[521].packet_type = "AXI_READ";
        traffic_data[521].size_bytes = 64;
        traffic_data[522].timestamp = 333;
        traffic_data[522].source_node = 2;
        traffic_data[522].dest_node = 8;
        traffic_data[522].packet_type = "AXI_READ";
        traffic_data[522].size_bytes = 64;
        traffic_data[523].timestamp = 334;
        traffic_data[523].source_node = 1;
        traffic_data[523].dest_node = 11;
        traffic_data[523].packet_type = "CHI_WRITE";
        traffic_data[523].size_bytes = 64;
        traffic_data[524].timestamp = 336;
        traffic_data[524].source_node = 6;
        traffic_data[524].dest_node = 12;
        traffic_data[524].packet_type = "AXI_READ";
        traffic_data[524].size_bytes = 64;
        traffic_data[525].timestamp = 336;
        traffic_data[525].source_node = 9;
        traffic_data[525].dest_node = 2;
        traffic_data[525].packet_type = "CHI_WRITE";
        traffic_data[525].size_bytes = 64;
        traffic_data[526].timestamp = 337;
        traffic_data[526].source_node = 9;
        traffic_data[526].dest_node = 13;
        traffic_data[526].packet_type = "AXI_READ";
        traffic_data[526].size_bytes = 64;
        traffic_data[527].timestamp = 338;
        traffic_data[527].source_node = 0;
        traffic_data[527].dest_node = 3;
        traffic_data[527].packet_type = "CHI_READ";
        traffic_data[527].size_bytes = 64;
        traffic_data[528].timestamp = 338;
        traffic_data[528].source_node = 14;
        traffic_data[528].dest_node = 4;
        traffic_data[528].packet_type = "CHI_WRITE";
        traffic_data[528].size_bytes = 64;
        traffic_data[529].timestamp = 339;
        traffic_data[529].source_node = 4;
        traffic_data[529].dest_node = 10;
        traffic_data[529].packet_type = "AXI_READ";
        traffic_data[529].size_bytes = 64;
        traffic_data[530].timestamp = 339;
        traffic_data[530].source_node = 15;
        traffic_data[530].dest_node = 3;
        traffic_data[530].packet_type = "AXI_WRITE";
        traffic_data[530].size_bytes = 64;
        traffic_data[531].timestamp = 340;
        traffic_data[531].source_node = 2;
        traffic_data[531].dest_node = 12;
        traffic_data[531].packet_type = "AXI_READ";
        traffic_data[531].size_bytes = 64;
        traffic_data[532].timestamp = 340;
        traffic_data[532].source_node = 7;
        traffic_data[532].dest_node = 11;
        traffic_data[532].packet_type = "CHI_WRITE";
        traffic_data[532].size_bytes = 64;
        traffic_data[533].timestamp = 342;
        traffic_data[533].source_node = 1;
        traffic_data[533].dest_node = 10;
        traffic_data[533].packet_type = "CHI_WRITE";
        traffic_data[533].size_bytes = 64;
        traffic_data[534].timestamp = 342;
        traffic_data[534].source_node = 13;
        traffic_data[534].dest_node = 14;
        traffic_data[534].packet_type = "CHI_READ";
        traffic_data[534].size_bytes = 64;
        traffic_data[535].timestamp = 344;
        traffic_data[535].source_node = 6;
        traffic_data[535].dest_node = 3;
        traffic_data[535].packet_type = "CHI_READ";
        traffic_data[535].size_bytes = 64;
        traffic_data[536].timestamp = 345;
        traffic_data[536].source_node = 8;
        traffic_data[536].dest_node = 13;
        traffic_data[536].packet_type = "CHI_READ";
        traffic_data[536].size_bytes = 64;
        traffic_data[537].timestamp = 345;
        traffic_data[537].source_node = 13;
        traffic_data[537].dest_node = 2;
        traffic_data[537].packet_type = "CHI_READ";
        traffic_data[537].size_bytes = 64;
        traffic_data[538].timestamp = 346;
        traffic_data[538].source_node = 6;
        traffic_data[538].dest_node = 14;
        traffic_data[538].packet_type = "AXI_READ";
        traffic_data[538].size_bytes = 64;
        traffic_data[539].timestamp = 346;
        traffic_data[539].source_node = 9;
        traffic_data[539].dest_node = 6;
        traffic_data[539].packet_type = "CHI_READ";
        traffic_data[539].size_bytes = 64;
        traffic_data[540].timestamp = 347;
        traffic_data[540].source_node = 8;
        traffic_data[540].dest_node = 10;
        traffic_data[540].packet_type = "AXI_READ";
        traffic_data[540].size_bytes = 64;
        traffic_data[541].timestamp = 348;
        traffic_data[541].source_node = 6;
        traffic_data[541].dest_node = 9;
        traffic_data[541].packet_type = "CHI_READ";
        traffic_data[541].size_bytes = 64;
        traffic_data[542].timestamp = 349;
        traffic_data[542].source_node = 4;
        traffic_data[542].dest_node = 12;
        traffic_data[542].packet_type = "AXI_READ";
        traffic_data[542].size_bytes = 64;
        traffic_data[543].timestamp = 350;
        traffic_data[543].source_node = 5;
        traffic_data[543].dest_node = 14;
        traffic_data[543].packet_type = "AXI_WRITE";
        traffic_data[543].size_bytes = 64;
        traffic_data[544].timestamp = 350;
        traffic_data[544].source_node = 15;
        traffic_data[544].dest_node = 12;
        traffic_data[544].packet_type = "CHI_WRITE";
        traffic_data[544].size_bytes = 64;
        traffic_data[545].timestamp = 351;
        traffic_data[545].source_node = 14;
        traffic_data[545].dest_node = 0;
        traffic_data[545].packet_type = "AXI_WRITE";
        traffic_data[545].size_bytes = 64;
        traffic_data[546].timestamp = 352;
        traffic_data[546].source_node = 5;
        traffic_data[546].dest_node = 2;
        traffic_data[546].packet_type = "AXI_WRITE";
        traffic_data[546].size_bytes = 64;
        traffic_data[547].timestamp = 354;
        traffic_data[547].source_node = 7;
        traffic_data[547].dest_node = 5;
        traffic_data[547].packet_type = "AXI_WRITE";
        traffic_data[547].size_bytes = 64;
        traffic_data[548].timestamp = 356;
        traffic_data[548].source_node = 6;
        traffic_data[548].dest_node = 2;
        traffic_data[548].packet_type = "CHI_READ";
        traffic_data[548].size_bytes = 64;
        traffic_data[549].timestamp = 356;
        traffic_data[549].source_node = 13;
        traffic_data[549].dest_node = 8;
        traffic_data[549].packet_type = "AXI_READ";
        traffic_data[549].size_bytes = 64;
        traffic_data[550].timestamp = 356;
        traffic_data[550].source_node = 14;
        traffic_data[550].dest_node = 15;
        traffic_data[550].packet_type = "AXI_WRITE";
        traffic_data[550].size_bytes = 64;
        traffic_data[551].timestamp = 357;
        traffic_data[551].source_node = 6;
        traffic_data[551].dest_node = 9;
        traffic_data[551].packet_type = "CHI_WRITE";
        traffic_data[551].size_bytes = 64;
        traffic_data[552].timestamp = 358;
        traffic_data[552].source_node = 6;
        traffic_data[552].dest_node = 2;
        traffic_data[552].packet_type = "CHI_WRITE";
        traffic_data[552].size_bytes = 64;
        traffic_data[553].timestamp = 359;
        traffic_data[553].source_node = 9;
        traffic_data[553].dest_node = 2;
        traffic_data[553].packet_type = "AXI_READ";
        traffic_data[553].size_bytes = 64;
        traffic_data[554].timestamp = 359;
        traffic_data[554].source_node = 11;
        traffic_data[554].dest_node = 4;
        traffic_data[554].packet_type = "AXI_WRITE";
        traffic_data[554].size_bytes = 64;
        traffic_data[555].timestamp = 360;
        traffic_data[555].source_node = 0;
        traffic_data[555].dest_node = 6;
        traffic_data[555].packet_type = "CHI_WRITE";
        traffic_data[555].size_bytes = 64;
        traffic_data[556].timestamp = 360;
        traffic_data[556].source_node = 15;
        traffic_data[556].dest_node = 12;
        traffic_data[556].packet_type = "AXI_WRITE";
        traffic_data[556].size_bytes = 64;
        traffic_data[557].timestamp = 361;
        traffic_data[557].source_node = 1;
        traffic_data[557].dest_node = 13;
        traffic_data[557].packet_type = "CHI_WRITE";
        traffic_data[557].size_bytes = 64;
        traffic_data[558].timestamp = 361;
        traffic_data[558].source_node = 4;
        traffic_data[558].dest_node = 11;
        traffic_data[558].packet_type = "AXI_READ";
        traffic_data[558].size_bytes = 64;
        traffic_data[559].timestamp = 361;
        traffic_data[559].source_node = 10;
        traffic_data[559].dest_node = 14;
        traffic_data[559].packet_type = "CHI_WRITE";
        traffic_data[559].size_bytes = 64;
        traffic_data[560].timestamp = 361;
        traffic_data[560].source_node = 14;
        traffic_data[560].dest_node = 0;
        traffic_data[560].packet_type = "CHI_WRITE";
        traffic_data[560].size_bytes = 64;
        traffic_data[561].timestamp = 362;
        traffic_data[561].source_node = 5;
        traffic_data[561].dest_node = 11;
        traffic_data[561].packet_type = "CHI_READ";
        traffic_data[561].size_bytes = 64;
        traffic_data[562].timestamp = 362;
        traffic_data[562].source_node = 7;
        traffic_data[562].dest_node = 1;
        traffic_data[562].packet_type = "CHI_WRITE";
        traffic_data[562].size_bytes = 64;
        traffic_data[563].timestamp = 362;
        traffic_data[563].source_node = 8;
        traffic_data[563].dest_node = 4;
        traffic_data[563].packet_type = "AXI_WRITE";
        traffic_data[563].size_bytes = 64;
        traffic_data[564].timestamp = 362;
        traffic_data[564].source_node = 12;
        traffic_data[564].dest_node = 3;
        traffic_data[564].packet_type = "AXI_WRITE";
        traffic_data[564].size_bytes = 64;
        traffic_data[565].timestamp = 363;
        traffic_data[565].source_node = 9;
        traffic_data[565].dest_node = 5;
        traffic_data[565].packet_type = "AXI_WRITE";
        traffic_data[565].size_bytes = 64;
        traffic_data[566].timestamp = 364;
        traffic_data[566].source_node = 4;
        traffic_data[566].dest_node = 6;
        traffic_data[566].packet_type = "CHI_WRITE";
        traffic_data[566].size_bytes = 64;
        traffic_data[567].timestamp = 364;
        traffic_data[567].source_node = 11;
        traffic_data[567].dest_node = 7;
        traffic_data[567].packet_type = "CHI_WRITE";
        traffic_data[567].size_bytes = 64;
        traffic_data[568].timestamp = 364;
        traffic_data[568].source_node = 12;
        traffic_data[568].dest_node = 13;
        traffic_data[568].packet_type = "CHI_WRITE";
        traffic_data[568].size_bytes = 64;
        traffic_data[569].timestamp = 365;
        traffic_data[569].source_node = 15;
        traffic_data[569].dest_node = 11;
        traffic_data[569].packet_type = "CHI_WRITE";
        traffic_data[569].size_bytes = 64;
        traffic_data[570].timestamp = 366;
        traffic_data[570].source_node = 3;
        traffic_data[570].dest_node = 15;
        traffic_data[570].packet_type = "CHI_READ";
        traffic_data[570].size_bytes = 64;
        traffic_data[571].timestamp = 366;
        traffic_data[571].source_node = 13;
        traffic_data[571].dest_node = 9;
        traffic_data[571].packet_type = "CHI_READ";
        traffic_data[571].size_bytes = 64;
        traffic_data[572].timestamp = 367;
        traffic_data[572].source_node = 1;
        traffic_data[572].dest_node = 2;
        traffic_data[572].packet_type = "AXI_READ";
        traffic_data[572].size_bytes = 64;
        traffic_data[573].timestamp = 368;
        traffic_data[573].source_node = 1;
        traffic_data[573].dest_node = 2;
        traffic_data[573].packet_type = "AXI_READ";
        traffic_data[573].size_bytes = 64;
        traffic_data[574].timestamp = 368;
        traffic_data[574].source_node = 4;
        traffic_data[574].dest_node = 8;
        traffic_data[574].packet_type = "AXI_WRITE";
        traffic_data[574].size_bytes = 64;
        traffic_data[575].timestamp = 368;
        traffic_data[575].source_node = 13;
        traffic_data[575].dest_node = 2;
        traffic_data[575].packet_type = "AXI_WRITE";
        traffic_data[575].size_bytes = 64;
        traffic_data[576].timestamp = 369;
        traffic_data[576].source_node = 1;
        traffic_data[576].dest_node = 8;
        traffic_data[576].packet_type = "AXI_WRITE";
        traffic_data[576].size_bytes = 64;
        traffic_data[577].timestamp = 369;
        traffic_data[577].source_node = 5;
        traffic_data[577].dest_node = 0;
        traffic_data[577].packet_type = "AXI_READ";
        traffic_data[577].size_bytes = 64;
        traffic_data[578].timestamp = 370;
        traffic_data[578].source_node = 9;
        traffic_data[578].dest_node = 15;
        traffic_data[578].packet_type = "CHI_WRITE";
        traffic_data[578].size_bytes = 64;
        traffic_data[579].timestamp = 372;
        traffic_data[579].source_node = 7;
        traffic_data[579].dest_node = 8;
        traffic_data[579].packet_type = "AXI_WRITE";
        traffic_data[579].size_bytes = 64;
        traffic_data[580].timestamp = 374;
        traffic_data[580].source_node = 7;
        traffic_data[580].dest_node = 8;
        traffic_data[580].packet_type = "CHI_WRITE";
        traffic_data[580].size_bytes = 64;
        traffic_data[581].timestamp = 376;
        traffic_data[581].source_node = 1;
        traffic_data[581].dest_node = 14;
        traffic_data[581].packet_type = "CHI_WRITE";
        traffic_data[581].size_bytes = 64;
        traffic_data[582].timestamp = 376;
        traffic_data[582].source_node = 4;
        traffic_data[582].dest_node = 6;
        traffic_data[582].packet_type = "CHI_WRITE";
        traffic_data[582].size_bytes = 64;
        traffic_data[583].timestamp = 377;
        traffic_data[583].source_node = 2;
        traffic_data[583].dest_node = 3;
        traffic_data[583].packet_type = "AXI_READ";
        traffic_data[583].size_bytes = 64;
        traffic_data[584].timestamp = 377;
        traffic_data[584].source_node = 5;
        traffic_data[584].dest_node = 6;
        traffic_data[584].packet_type = "CHI_READ";
        traffic_data[584].size_bytes = 64;
        traffic_data[585].timestamp = 377;
        traffic_data[585].source_node = 10;
        traffic_data[585].dest_node = 15;
        traffic_data[585].packet_type = "AXI_WRITE";
        traffic_data[585].size_bytes = 64;
        traffic_data[586].timestamp = 377;
        traffic_data[586].source_node = 12;
        traffic_data[586].dest_node = 10;
        traffic_data[586].packet_type = "CHI_READ";
        traffic_data[586].size_bytes = 64;
        traffic_data[587].timestamp = 379;
        traffic_data[587].source_node = 3;
        traffic_data[587].dest_node = 9;
        traffic_data[587].packet_type = "CHI_READ";
        traffic_data[587].size_bytes = 64;
        traffic_data[588].timestamp = 379;
        traffic_data[588].source_node = 14;
        traffic_data[588].dest_node = 15;
        traffic_data[588].packet_type = "CHI_READ";
        traffic_data[588].size_bytes = 64;
        traffic_data[589].timestamp = 380;
        traffic_data[589].source_node = 4;
        traffic_data[589].dest_node = 6;
        traffic_data[589].packet_type = "CHI_READ";
        traffic_data[589].size_bytes = 64;
        traffic_data[590].timestamp = 380;
        traffic_data[590].source_node = 7;
        traffic_data[590].dest_node = 11;
        traffic_data[590].packet_type = "AXI_READ";
        traffic_data[590].size_bytes = 64;
        traffic_data[591].timestamp = 380;
        traffic_data[591].source_node = 10;
        traffic_data[591].dest_node = 5;
        traffic_data[591].packet_type = "AXI_WRITE";
        traffic_data[591].size_bytes = 64;
        traffic_data[592].timestamp = 381;
        traffic_data[592].source_node = 14;
        traffic_data[592].dest_node = 11;
        traffic_data[592].packet_type = "CHI_WRITE";
        traffic_data[592].size_bytes = 64;
        traffic_data[593].timestamp = 382;
        traffic_data[593].source_node = 0;
        traffic_data[593].dest_node = 1;
        traffic_data[593].packet_type = "CHI_WRITE";
        traffic_data[593].size_bytes = 64;
        traffic_data[594].timestamp = 384;
        traffic_data[594].source_node = 2;
        traffic_data[594].dest_node = 3;
        traffic_data[594].packet_type = "AXI_READ";
        traffic_data[594].size_bytes = 64;
        traffic_data[595].timestamp = 384;
        traffic_data[595].source_node = 10;
        traffic_data[595].dest_node = 15;
        traffic_data[595].packet_type = "CHI_READ";
        traffic_data[595].size_bytes = 64;
        traffic_data[596].timestamp = 387;
        traffic_data[596].source_node = 6;
        traffic_data[596].dest_node = 10;
        traffic_data[596].packet_type = "AXI_WRITE";
        traffic_data[596].size_bytes = 64;
        traffic_data[597].timestamp = 387;
        traffic_data[597].source_node = 9;
        traffic_data[597].dest_node = 11;
        traffic_data[597].packet_type = "AXI_WRITE";
        traffic_data[597].size_bytes = 64;
        traffic_data[598].timestamp = 388;
        traffic_data[598].source_node = 0;
        traffic_data[598].dest_node = 9;
        traffic_data[598].packet_type = "CHI_READ";
        traffic_data[598].size_bytes = 64;
        traffic_data[599].timestamp = 388;
        traffic_data[599].source_node = 2;
        traffic_data[599].dest_node = 14;
        traffic_data[599].packet_type = "AXI_READ";
        traffic_data[599].size_bytes = 64;
        traffic_data[600].timestamp = 388;
        traffic_data[600].source_node = 5;
        traffic_data[600].dest_node = 9;
        traffic_data[600].packet_type = "CHI_READ";
        traffic_data[600].size_bytes = 64;
        traffic_data[601].timestamp = 388;
        traffic_data[601].source_node = 7;
        traffic_data[601].dest_node = 1;
        traffic_data[601].packet_type = "AXI_WRITE";
        traffic_data[601].size_bytes = 64;
        traffic_data[602].timestamp = 388;
        traffic_data[602].source_node = 14;
        traffic_data[602].dest_node = 5;
        traffic_data[602].packet_type = "AXI_WRITE";
        traffic_data[602].size_bytes = 64;
        traffic_data[603].timestamp = 388;
        traffic_data[603].source_node = 15;
        traffic_data[603].dest_node = 0;
        traffic_data[603].packet_type = "CHI_READ";
        traffic_data[603].size_bytes = 64;
        traffic_data[604].timestamp = 389;
        traffic_data[604].source_node = 14;
        traffic_data[604].dest_node = 7;
        traffic_data[604].packet_type = "CHI_WRITE";
        traffic_data[604].size_bytes = 64;
        traffic_data[605].timestamp = 389;
        traffic_data[605].source_node = 15;
        traffic_data[605].dest_node = 0;
        traffic_data[605].packet_type = "CHI_WRITE";
        traffic_data[605].size_bytes = 64;
        traffic_data[606].timestamp = 390;
        traffic_data[606].source_node = 2;
        traffic_data[606].dest_node = 9;
        traffic_data[606].packet_type = "AXI_READ";
        traffic_data[606].size_bytes = 64;
        traffic_data[607].timestamp = 390;
        traffic_data[607].source_node = 8;
        traffic_data[607].dest_node = 11;
        traffic_data[607].packet_type = "AXI_WRITE";
        traffic_data[607].size_bytes = 64;
        traffic_data[608].timestamp = 391;
        traffic_data[608].source_node = 1;
        traffic_data[608].dest_node = 14;
        traffic_data[608].packet_type = "CHI_WRITE";
        traffic_data[608].size_bytes = 64;
        traffic_data[609].timestamp = 391;
        traffic_data[609].source_node = 6;
        traffic_data[609].dest_node = 15;
        traffic_data[609].packet_type = "CHI_WRITE";
        traffic_data[609].size_bytes = 64;
        traffic_data[610].timestamp = 392;
        traffic_data[610].source_node = 1;
        traffic_data[610].dest_node = 2;
        traffic_data[610].packet_type = "CHI_WRITE";
        traffic_data[610].size_bytes = 64;
        traffic_data[611].timestamp = 393;
        traffic_data[611].source_node = 9;
        traffic_data[611].dest_node = 0;
        traffic_data[611].packet_type = "AXI_WRITE";
        traffic_data[611].size_bytes = 64;
        traffic_data[612].timestamp = 394;
        traffic_data[612].source_node = 1;
        traffic_data[612].dest_node = 0;
        traffic_data[612].packet_type = "CHI_WRITE";
        traffic_data[612].size_bytes = 64;
        traffic_data[613].timestamp = 394;
        traffic_data[613].source_node = 10;
        traffic_data[613].dest_node = 7;
        traffic_data[613].packet_type = "CHI_READ";
        traffic_data[613].size_bytes = 64;
        traffic_data[614].timestamp = 394;
        traffic_data[614].source_node = 14;
        traffic_data[614].dest_node = 4;
        traffic_data[614].packet_type = "CHI_READ";
        traffic_data[614].size_bytes = 64;
        traffic_data[615].timestamp = 395;
        traffic_data[615].source_node = 6;
        traffic_data[615].dest_node = 8;
        traffic_data[615].packet_type = "AXI_WRITE";
        traffic_data[615].size_bytes = 64;
        traffic_data[616].timestamp = 395;
        traffic_data[616].source_node = 7;
        traffic_data[616].dest_node = 14;
        traffic_data[616].packet_type = "CHI_WRITE";
        traffic_data[616].size_bytes = 64;
        traffic_data[617].timestamp = 396;
        traffic_data[617].source_node = 10;
        traffic_data[617].dest_node = 12;
        traffic_data[617].packet_type = "CHI_READ";
        traffic_data[617].size_bytes = 64;
        traffic_data[618].timestamp = 396;
        traffic_data[618].source_node = 13;
        traffic_data[618].dest_node = 6;
        traffic_data[618].packet_type = "AXI_READ";
        traffic_data[618].size_bytes = 64;
        traffic_data[619].timestamp = 397;
        traffic_data[619].source_node = 6;
        traffic_data[619].dest_node = 12;
        traffic_data[619].packet_type = "AXI_WRITE";
        traffic_data[619].size_bytes = 64;
        traffic_data[620].timestamp = 397;
        traffic_data[620].source_node = 7;
        traffic_data[620].dest_node = 15;
        traffic_data[620].packet_type = "CHI_WRITE";
        traffic_data[620].size_bytes = 64;
        traffic_data[621].timestamp = 398;
        traffic_data[621].source_node = 5;
        traffic_data[621].dest_node = 11;
        traffic_data[621].packet_type = "AXI_READ";
        traffic_data[621].size_bytes = 64;
        traffic_data[622].timestamp = 398;
        traffic_data[622].source_node = 6;
        traffic_data[622].dest_node = 7;
        traffic_data[622].packet_type = "AXI_READ";
        traffic_data[622].size_bytes = 64;
        traffic_data[623].timestamp = 398;
        traffic_data[623].source_node = 14;
        traffic_data[623].dest_node = 5;
        traffic_data[623].packet_type = "AXI_WRITE";
        traffic_data[623].size_bytes = 64;
        traffic_data[624].timestamp = 399;
        traffic_data[624].source_node = 5;
        traffic_data[624].dest_node = 0;
        traffic_data[624].packet_type = "AXI_READ";
        traffic_data[624].size_bytes = 64;
        traffic_data[625].timestamp = 399;
        traffic_data[625].source_node = 10;
        traffic_data[625].dest_node = 13;
        traffic_data[625].packet_type = "CHI_WRITE";
        traffic_data[625].size_bytes = 64;
        traffic_data[626].timestamp = 399;
        traffic_data[626].source_node = 11;
        traffic_data[626].dest_node = 9;
        traffic_data[626].packet_type = "CHI_WRITE";
        traffic_data[626].size_bytes = 64;
        traffic_data[627].timestamp = 399;
        traffic_data[627].source_node = 12;
        traffic_data[627].dest_node = 10;
        traffic_data[627].packet_type = "AXI_READ";
        traffic_data[627].size_bytes = 64;
        traffic_data[628].timestamp = 400;
        traffic_data[628].source_node = 0;
        traffic_data[628].dest_node = 13;
        traffic_data[628].packet_type = "CHI_WRITE";
        traffic_data[628].size_bytes = 64;
        traffic_data[629].timestamp = 400;
        traffic_data[629].source_node = 4;
        traffic_data[629].dest_node = 7;
        traffic_data[629].packet_type = "CHI_WRITE";
        traffic_data[629].size_bytes = 64;
        traffic_data[630].timestamp = 401;
        traffic_data[630].source_node = 0;
        traffic_data[630].dest_node = 13;
        traffic_data[630].packet_type = "AXI_WRITE";
        traffic_data[630].size_bytes = 64;
        traffic_data[631].timestamp = 401;
        traffic_data[631].source_node = 9;
        traffic_data[631].dest_node = 2;
        traffic_data[631].packet_type = "CHI_READ";
        traffic_data[631].size_bytes = 64;
        traffic_data[632].timestamp = 402;
        traffic_data[632].source_node = 11;
        traffic_data[632].dest_node = 5;
        traffic_data[632].packet_type = "AXI_WRITE";
        traffic_data[632].size_bytes = 64;
        traffic_data[633].timestamp = 402;
        traffic_data[633].source_node = 15;
        traffic_data[633].dest_node = 3;
        traffic_data[633].packet_type = "CHI_WRITE";
        traffic_data[633].size_bytes = 64;
        traffic_data[634].timestamp = 403;
        traffic_data[634].source_node = 11;
        traffic_data[634].dest_node = 3;
        traffic_data[634].packet_type = "AXI_READ";
        traffic_data[634].size_bytes = 64;
        traffic_data[635].timestamp = 404;
        traffic_data[635].source_node = 7;
        traffic_data[635].dest_node = 0;
        traffic_data[635].packet_type = "AXI_READ";
        traffic_data[635].size_bytes = 64;
        traffic_data[636].timestamp = 409;
        traffic_data[636].source_node = 14;
        traffic_data[636].dest_node = 12;
        traffic_data[636].packet_type = "AXI_READ";
        traffic_data[636].size_bytes = 64;
        traffic_data[637].timestamp = 410;
        traffic_data[637].source_node = 2;
        traffic_data[637].dest_node = 9;
        traffic_data[637].packet_type = "CHI_READ";
        traffic_data[637].size_bytes = 64;
        traffic_data[638].timestamp = 410;
        traffic_data[638].source_node = 13;
        traffic_data[638].dest_node = 14;
        traffic_data[638].packet_type = "AXI_READ";
        traffic_data[638].size_bytes = 64;
        traffic_data[639].timestamp = 411;
        traffic_data[639].source_node = 0;
        traffic_data[639].dest_node = 2;
        traffic_data[639].packet_type = "CHI_READ";
        traffic_data[639].size_bytes = 64;
        traffic_data[640].timestamp = 411;
        traffic_data[640].source_node = 1;
        traffic_data[640].dest_node = 4;
        traffic_data[640].packet_type = "CHI_READ";
        traffic_data[640].size_bytes = 64;
        traffic_data[641].timestamp = 411;
        traffic_data[641].source_node = 14;
        traffic_data[641].dest_node = 4;
        traffic_data[641].packet_type = "CHI_READ";
        traffic_data[641].size_bytes = 64;
        traffic_data[642].timestamp = 413;
        traffic_data[642].source_node = 14;
        traffic_data[642].dest_node = 12;
        traffic_data[642].packet_type = "CHI_READ";
        traffic_data[642].size_bytes = 64;
        traffic_data[643].timestamp = 414;
        traffic_data[643].source_node = 6;
        traffic_data[643].dest_node = 13;
        traffic_data[643].packet_type = "AXI_READ";
        traffic_data[643].size_bytes = 64;
        traffic_data[644].timestamp = 415;
        traffic_data[644].source_node = 8;
        traffic_data[644].dest_node = 1;
        traffic_data[644].packet_type = "AXI_WRITE";
        traffic_data[644].size_bytes = 64;
        traffic_data[645].timestamp = 415;
        traffic_data[645].source_node = 9;
        traffic_data[645].dest_node = 12;
        traffic_data[645].packet_type = "CHI_WRITE";
        traffic_data[645].size_bytes = 64;
        traffic_data[646].timestamp = 415;
        traffic_data[646].source_node = 10;
        traffic_data[646].dest_node = 3;
        traffic_data[646].packet_type = "AXI_READ";
        traffic_data[646].size_bytes = 64;
        traffic_data[647].timestamp = 416;
        traffic_data[647].source_node = 2;
        traffic_data[647].dest_node = 6;
        traffic_data[647].packet_type = "CHI_WRITE";
        traffic_data[647].size_bytes = 64;
        traffic_data[648].timestamp = 417;
        traffic_data[648].source_node = 15;
        traffic_data[648].dest_node = 1;
        traffic_data[648].packet_type = "CHI_READ";
        traffic_data[648].size_bytes = 64;
        traffic_data[649].timestamp = 418;
        traffic_data[649].source_node = 15;
        traffic_data[649].dest_node = 11;
        traffic_data[649].packet_type = "AXI_READ";
        traffic_data[649].size_bytes = 64;
        traffic_data[650].timestamp = 419;
        traffic_data[650].source_node = 13;
        traffic_data[650].dest_node = 1;
        traffic_data[650].packet_type = "CHI_READ";
        traffic_data[650].size_bytes = 64;
        traffic_data[651].timestamp = 420;
        traffic_data[651].source_node = 1;
        traffic_data[651].dest_node = 0;
        traffic_data[651].packet_type = "AXI_READ";
        traffic_data[651].size_bytes = 64;
        traffic_data[652].timestamp = 420;
        traffic_data[652].source_node = 8;
        traffic_data[652].dest_node = 4;
        traffic_data[652].packet_type = "AXI_READ";
        traffic_data[652].size_bytes = 64;
        traffic_data[653].timestamp = 420;
        traffic_data[653].source_node = 14;
        traffic_data[653].dest_node = 10;
        traffic_data[653].packet_type = "AXI_WRITE";
        traffic_data[653].size_bytes = 64;
        traffic_data[654].timestamp = 421;
        traffic_data[654].source_node = 11;
        traffic_data[654].dest_node = 4;
        traffic_data[654].packet_type = "AXI_WRITE";
        traffic_data[654].size_bytes = 64;
        traffic_data[655].timestamp = 422;
        traffic_data[655].source_node = 2;
        traffic_data[655].dest_node = 11;
        traffic_data[655].packet_type = "AXI_READ";
        traffic_data[655].size_bytes = 64;
        traffic_data[656].timestamp = 422;
        traffic_data[656].source_node = 5;
        traffic_data[656].dest_node = 0;
        traffic_data[656].packet_type = "AXI_READ";
        traffic_data[656].size_bytes = 64;
        traffic_data[657].timestamp = 422;
        traffic_data[657].source_node = 11;
        traffic_data[657].dest_node = 6;
        traffic_data[657].packet_type = "AXI_READ";
        traffic_data[657].size_bytes = 64;
        traffic_data[658].timestamp = 424;
        traffic_data[658].source_node = 6;
        traffic_data[658].dest_node = 14;
        traffic_data[658].packet_type = "CHI_READ";
        traffic_data[658].size_bytes = 64;
        traffic_data[659].timestamp = 424;
        traffic_data[659].source_node = 9;
        traffic_data[659].dest_node = 3;
        traffic_data[659].packet_type = "CHI_WRITE";
        traffic_data[659].size_bytes = 64;
        traffic_data[660].timestamp = 426;
        traffic_data[660].source_node = 14;
        traffic_data[660].dest_node = 5;
        traffic_data[660].packet_type = "CHI_WRITE";
        traffic_data[660].size_bytes = 64;
        traffic_data[661].timestamp = 427;
        traffic_data[661].source_node = 2;
        traffic_data[661].dest_node = 15;
        traffic_data[661].packet_type = "CHI_WRITE";
        traffic_data[661].size_bytes = 64;
        traffic_data[662].timestamp = 427;
        traffic_data[662].source_node = 12;
        traffic_data[662].dest_node = 14;
        traffic_data[662].packet_type = "CHI_READ";
        traffic_data[662].size_bytes = 64;
        traffic_data[663].timestamp = 427;
        traffic_data[663].source_node = 15;
        traffic_data[663].dest_node = 14;
        traffic_data[663].packet_type = "AXI_WRITE";
        traffic_data[663].size_bytes = 64;
        traffic_data[664].timestamp = 428;
        traffic_data[664].source_node = 7;
        traffic_data[664].dest_node = 8;
        traffic_data[664].packet_type = "AXI_READ";
        traffic_data[664].size_bytes = 64;
        traffic_data[665].timestamp = 428;
        traffic_data[665].source_node = 9;
        traffic_data[665].dest_node = 2;
        traffic_data[665].packet_type = "AXI_WRITE";
        traffic_data[665].size_bytes = 64;
        traffic_data[666].timestamp = 430;
        traffic_data[666].source_node = 8;
        traffic_data[666].dest_node = 15;
        traffic_data[666].packet_type = "CHI_READ";
        traffic_data[666].size_bytes = 64;
        traffic_data[667].timestamp = 431;
        traffic_data[667].source_node = 1;
        traffic_data[667].dest_node = 3;
        traffic_data[667].packet_type = "CHI_WRITE";
        traffic_data[667].size_bytes = 64;
        traffic_data[668].timestamp = 431;
        traffic_data[668].source_node = 4;
        traffic_data[668].dest_node = 14;
        traffic_data[668].packet_type = "CHI_READ";
        traffic_data[668].size_bytes = 64;
        traffic_data[669].timestamp = 431;
        traffic_data[669].source_node = 14;
        traffic_data[669].dest_node = 15;
        traffic_data[669].packet_type = "AXI_READ";
        traffic_data[669].size_bytes = 64;
        traffic_data[670].timestamp = 432;
        traffic_data[670].source_node = 14;
        traffic_data[670].dest_node = 13;
        traffic_data[670].packet_type = "CHI_READ";
        traffic_data[670].size_bytes = 64;
        traffic_data[671].timestamp = 433;
        traffic_data[671].source_node = 10;
        traffic_data[671].dest_node = 13;
        traffic_data[671].packet_type = "AXI_READ";
        traffic_data[671].size_bytes = 64;
        traffic_data[672].timestamp = 434;
        traffic_data[672].source_node = 13;
        traffic_data[672].dest_node = 10;
        traffic_data[672].packet_type = "CHI_READ";
        traffic_data[672].size_bytes = 64;
        traffic_data[673].timestamp = 435;
        traffic_data[673].source_node = 3;
        traffic_data[673].dest_node = 2;
        traffic_data[673].packet_type = "CHI_WRITE";
        traffic_data[673].size_bytes = 64;
        traffic_data[674].timestamp = 435;
        traffic_data[674].source_node = 4;
        traffic_data[674].dest_node = 1;
        traffic_data[674].packet_type = "CHI_WRITE";
        traffic_data[674].size_bytes = 64;
        traffic_data[675].timestamp = 436;
        traffic_data[675].source_node = 1;
        traffic_data[675].dest_node = 3;
        traffic_data[675].packet_type = "AXI_WRITE";
        traffic_data[675].size_bytes = 64;
        traffic_data[676].timestamp = 437;
        traffic_data[676].source_node = 1;
        traffic_data[676].dest_node = 13;
        traffic_data[676].packet_type = "AXI_READ";
        traffic_data[676].size_bytes = 64;
        traffic_data[677].timestamp = 437;
        traffic_data[677].source_node = 4;
        traffic_data[677].dest_node = 3;
        traffic_data[677].packet_type = "AXI_READ";
        traffic_data[677].size_bytes = 64;
        traffic_data[678].timestamp = 438;
        traffic_data[678].source_node = 7;
        traffic_data[678].dest_node = 14;
        traffic_data[678].packet_type = "CHI_WRITE";
        traffic_data[678].size_bytes = 64;
        traffic_data[679].timestamp = 439;
        traffic_data[679].source_node = 9;
        traffic_data[679].dest_node = 5;
        traffic_data[679].packet_type = "AXI_READ";
        traffic_data[679].size_bytes = 64;
        traffic_data[680].timestamp = 440;
        traffic_data[680].source_node = 15;
        traffic_data[680].dest_node = 7;
        traffic_data[680].packet_type = "AXI_READ";
        traffic_data[680].size_bytes = 64;
        traffic_data[681].timestamp = 441;
        traffic_data[681].source_node = 12;
        traffic_data[681].dest_node = 6;
        traffic_data[681].packet_type = "AXI_READ";
        traffic_data[681].size_bytes = 64;
        traffic_data[682].timestamp = 442;
        traffic_data[682].source_node = 9;
        traffic_data[682].dest_node = 12;
        traffic_data[682].packet_type = "CHI_READ";
        traffic_data[682].size_bytes = 64;
        traffic_data[683].timestamp = 443;
        traffic_data[683].source_node = 9;
        traffic_data[683].dest_node = 1;
        traffic_data[683].packet_type = "CHI_READ";
        traffic_data[683].size_bytes = 64;
        traffic_data[684].timestamp = 444;
        traffic_data[684].source_node = 2;
        traffic_data[684].dest_node = 0;
        traffic_data[684].packet_type = "AXI_WRITE";
        traffic_data[684].size_bytes = 64;
        traffic_data[685].timestamp = 446;
        traffic_data[685].source_node = 11;
        traffic_data[685].dest_node = 14;
        traffic_data[685].packet_type = "AXI_WRITE";
        traffic_data[685].size_bytes = 64;
        traffic_data[686].timestamp = 447;
        traffic_data[686].source_node = 2;
        traffic_data[686].dest_node = 7;
        traffic_data[686].packet_type = "CHI_READ";
        traffic_data[686].size_bytes = 64;
        traffic_data[687].timestamp = 447;
        traffic_data[687].source_node = 7;
        traffic_data[687].dest_node = 12;
        traffic_data[687].packet_type = "CHI_READ";
        traffic_data[687].size_bytes = 64;
        traffic_data[688].timestamp = 447;
        traffic_data[688].source_node = 12;
        traffic_data[688].dest_node = 5;
        traffic_data[688].packet_type = "AXI_READ";
        traffic_data[688].size_bytes = 64;
        traffic_data[689].timestamp = 448;
        traffic_data[689].source_node = 8;
        traffic_data[689].dest_node = 12;
        traffic_data[689].packet_type = "AXI_READ";
        traffic_data[689].size_bytes = 64;
        traffic_data[690].timestamp = 449;
        traffic_data[690].source_node = 0;
        traffic_data[690].dest_node = 8;
        traffic_data[690].packet_type = "AXI_WRITE";
        traffic_data[690].size_bytes = 64;
        traffic_data[691].timestamp = 450;
        traffic_data[691].source_node = 2;
        traffic_data[691].dest_node = 8;
        traffic_data[691].packet_type = "CHI_WRITE";
        traffic_data[691].size_bytes = 64;
        traffic_data[692].timestamp = 450;
        traffic_data[692].source_node = 7;
        traffic_data[692].dest_node = 8;
        traffic_data[692].packet_type = "AXI_WRITE";
        traffic_data[692].size_bytes = 64;
        traffic_data[693].timestamp = 450;
        traffic_data[693].source_node = 8;
        traffic_data[693].dest_node = 10;
        traffic_data[693].packet_type = "CHI_WRITE";
        traffic_data[693].size_bytes = 64;
        traffic_data[694].timestamp = 451;
        traffic_data[694].source_node = 1;
        traffic_data[694].dest_node = 2;
        traffic_data[694].packet_type = "AXI_WRITE";
        traffic_data[694].size_bytes = 64;
        traffic_data[695].timestamp = 451;
        traffic_data[695].source_node = 8;
        traffic_data[695].dest_node = 14;
        traffic_data[695].packet_type = "AXI_READ";
        traffic_data[695].size_bytes = 64;
        traffic_data[696].timestamp = 451;
        traffic_data[696].source_node = 15;
        traffic_data[696].dest_node = 7;
        traffic_data[696].packet_type = "CHI_READ";
        traffic_data[696].size_bytes = 64;
        traffic_data[697].timestamp = 452;
        traffic_data[697].source_node = 6;
        traffic_data[697].dest_node = 1;
        traffic_data[697].packet_type = "CHI_READ";
        traffic_data[697].size_bytes = 64;
        traffic_data[698].timestamp = 452;
        traffic_data[698].source_node = 11;
        traffic_data[698].dest_node = 4;
        traffic_data[698].packet_type = "AXI_READ";
        traffic_data[698].size_bytes = 64;
        traffic_data[699].timestamp = 453;
        traffic_data[699].source_node = 8;
        traffic_data[699].dest_node = 14;
        traffic_data[699].packet_type = "AXI_READ";
        traffic_data[699].size_bytes = 64;
        traffic_data[700].timestamp = 454;
        traffic_data[700].source_node = 3;
        traffic_data[700].dest_node = 5;
        traffic_data[700].packet_type = "CHI_READ";
        traffic_data[700].size_bytes = 64;
        traffic_data[701].timestamp = 454;
        traffic_data[701].source_node = 7;
        traffic_data[701].dest_node = 4;
        traffic_data[701].packet_type = "CHI_WRITE";
        traffic_data[701].size_bytes = 64;
        traffic_data[702].timestamp = 455;
        traffic_data[702].source_node = 15;
        traffic_data[702].dest_node = 14;
        traffic_data[702].packet_type = "CHI_READ";
        traffic_data[702].size_bytes = 64;
        traffic_data[703].timestamp = 456;
        traffic_data[703].source_node = 4;
        traffic_data[703].dest_node = 3;
        traffic_data[703].packet_type = "CHI_WRITE";
        traffic_data[703].size_bytes = 64;
        traffic_data[704].timestamp = 456;
        traffic_data[704].source_node = 12;
        traffic_data[704].dest_node = 5;
        traffic_data[704].packet_type = "CHI_READ";
        traffic_data[704].size_bytes = 64;
        traffic_data[705].timestamp = 457;
        traffic_data[705].source_node = 11;
        traffic_data[705].dest_node = 8;
        traffic_data[705].packet_type = "AXI_WRITE";
        traffic_data[705].size_bytes = 64;
        traffic_data[706].timestamp = 459;
        traffic_data[706].source_node = 1;
        traffic_data[706].dest_node = 5;
        traffic_data[706].packet_type = "CHI_WRITE";
        traffic_data[706].size_bytes = 64;
        traffic_data[707].timestamp = 459;
        traffic_data[707].source_node = 5;
        traffic_data[707].dest_node = 3;
        traffic_data[707].packet_type = "AXI_READ";
        traffic_data[707].size_bytes = 64;
        traffic_data[708].timestamp = 459;
        traffic_data[708].source_node = 7;
        traffic_data[708].dest_node = 12;
        traffic_data[708].packet_type = "CHI_READ";
        traffic_data[708].size_bytes = 64;
        traffic_data[709].timestamp = 461;
        traffic_data[709].source_node = 8;
        traffic_data[709].dest_node = 14;
        traffic_data[709].packet_type = "AXI_WRITE";
        traffic_data[709].size_bytes = 64;
        traffic_data[710].timestamp = 462;
        traffic_data[710].source_node = 14;
        traffic_data[710].dest_node = 7;
        traffic_data[710].packet_type = "CHI_WRITE";
        traffic_data[710].size_bytes = 64;
        traffic_data[711].timestamp = 462;
        traffic_data[711].source_node = 15;
        traffic_data[711].dest_node = 0;
        traffic_data[711].packet_type = "CHI_WRITE";
        traffic_data[711].size_bytes = 64;
        traffic_data[712].timestamp = 463;
        traffic_data[712].source_node = 2;
        traffic_data[712].dest_node = 15;
        traffic_data[712].packet_type = "AXI_WRITE";
        traffic_data[712].size_bytes = 64;
        traffic_data[713].timestamp = 463;
        traffic_data[713].source_node = 4;
        traffic_data[713].dest_node = 7;
        traffic_data[713].packet_type = "CHI_WRITE";
        traffic_data[713].size_bytes = 64;
        traffic_data[714].timestamp = 463;
        traffic_data[714].source_node = 10;
        traffic_data[714].dest_node = 13;
        traffic_data[714].packet_type = "CHI_READ";
        traffic_data[714].size_bytes = 64;
        traffic_data[715].timestamp = 464;
        traffic_data[715].source_node = 11;
        traffic_data[715].dest_node = 6;
        traffic_data[715].packet_type = "CHI_WRITE";
        traffic_data[715].size_bytes = 64;
        traffic_data[716].timestamp = 466;
        traffic_data[716].source_node = 0;
        traffic_data[716].dest_node = 3;
        traffic_data[716].packet_type = "CHI_READ";
        traffic_data[716].size_bytes = 64;
        traffic_data[717].timestamp = 468;
        traffic_data[717].source_node = 0;
        traffic_data[717].dest_node = 4;
        traffic_data[717].packet_type = "AXI_WRITE";
        traffic_data[717].size_bytes = 64;
        traffic_data[718].timestamp = 468;
        traffic_data[718].source_node = 3;
        traffic_data[718].dest_node = 0;
        traffic_data[718].packet_type = "CHI_WRITE";
        traffic_data[718].size_bytes = 64;
        traffic_data[719].timestamp = 469;
        traffic_data[719].source_node = 2;
        traffic_data[719].dest_node = 0;
        traffic_data[719].packet_type = "AXI_READ";
        traffic_data[719].size_bytes = 64;
        traffic_data[720].timestamp = 469;
        traffic_data[720].source_node = 3;
        traffic_data[720].dest_node = 12;
        traffic_data[720].packet_type = "CHI_READ";
        traffic_data[720].size_bytes = 64;
        traffic_data[721].timestamp = 469;
        traffic_data[721].source_node = 12;
        traffic_data[721].dest_node = 0;
        traffic_data[721].packet_type = "AXI_WRITE";
        traffic_data[721].size_bytes = 64;
        traffic_data[722].timestamp = 471;
        traffic_data[722].source_node = 0;
        traffic_data[722].dest_node = 9;
        traffic_data[722].packet_type = "CHI_READ";
        traffic_data[722].size_bytes = 64;
        traffic_data[723].timestamp = 472;
        traffic_data[723].source_node = 11;
        traffic_data[723].dest_node = 12;
        traffic_data[723].packet_type = "AXI_WRITE";
        traffic_data[723].size_bytes = 64;
        traffic_data[724].timestamp = 474;
        traffic_data[724].source_node = 5;
        traffic_data[724].dest_node = 3;
        traffic_data[724].packet_type = "CHI_READ";
        traffic_data[724].size_bytes = 64;
        traffic_data[725].timestamp = 474;
        traffic_data[725].source_node = 6;
        traffic_data[725].dest_node = 2;
        traffic_data[725].packet_type = "CHI_READ";
        traffic_data[725].size_bytes = 64;
        traffic_data[726].timestamp = 474;
        traffic_data[726].source_node = 14;
        traffic_data[726].dest_node = 5;
        traffic_data[726].packet_type = "CHI_READ";
        traffic_data[726].size_bytes = 64;
        traffic_data[727].timestamp = 475;
        traffic_data[727].source_node = 8;
        traffic_data[727].dest_node = 5;
        traffic_data[727].packet_type = "AXI_WRITE";
        traffic_data[727].size_bytes = 64;
        traffic_data[728].timestamp = 475;
        traffic_data[728].source_node = 12;
        traffic_data[728].dest_node = 10;
        traffic_data[728].packet_type = "AXI_READ";
        traffic_data[728].size_bytes = 64;
        traffic_data[729].timestamp = 478;
        traffic_data[729].source_node = 4;
        traffic_data[729].dest_node = 1;
        traffic_data[729].packet_type = "CHI_WRITE";
        traffic_data[729].size_bytes = 64;
        traffic_data[730].timestamp = 478;
        traffic_data[730].source_node = 7;
        traffic_data[730].dest_node = 14;
        traffic_data[730].packet_type = "AXI_READ";
        traffic_data[730].size_bytes = 64;
        traffic_data[731].timestamp = 478;
        traffic_data[731].source_node = 14;
        traffic_data[731].dest_node = 12;
        traffic_data[731].packet_type = "AXI_READ";
        traffic_data[731].size_bytes = 64;
        traffic_data[732].timestamp = 479;
        traffic_data[732].source_node = 2;
        traffic_data[732].dest_node = 3;
        traffic_data[732].packet_type = "CHI_WRITE";
        traffic_data[732].size_bytes = 64;
        traffic_data[733].timestamp = 479;
        traffic_data[733].source_node = 12;
        traffic_data[733].dest_node = 0;
        traffic_data[733].packet_type = "AXI_READ";
        traffic_data[733].size_bytes = 64;
        traffic_data[734].timestamp = 480;
        traffic_data[734].source_node = 1;
        traffic_data[734].dest_node = 4;
        traffic_data[734].packet_type = "AXI_READ";
        traffic_data[734].size_bytes = 64;
        traffic_data[735].timestamp = 481;
        traffic_data[735].source_node = 0;
        traffic_data[735].dest_node = 6;
        traffic_data[735].packet_type = "AXI_READ";
        traffic_data[735].size_bytes = 64;
        traffic_data[736].timestamp = 481;
        traffic_data[736].source_node = 3;
        traffic_data[736].dest_node = 0;
        traffic_data[736].packet_type = "AXI_WRITE";
        traffic_data[736].size_bytes = 64;
        traffic_data[737].timestamp = 482;
        traffic_data[737].source_node = 3;
        traffic_data[737].dest_node = 0;
        traffic_data[737].packet_type = "AXI_WRITE";
        traffic_data[737].size_bytes = 64;
        traffic_data[738].timestamp = 484;
        traffic_data[738].source_node = 1;
        traffic_data[738].dest_node = 12;
        traffic_data[738].packet_type = "CHI_WRITE";
        traffic_data[738].size_bytes = 64;
        traffic_data[739].timestamp = 484;
        traffic_data[739].source_node = 6;
        traffic_data[739].dest_node = 5;
        traffic_data[739].packet_type = "AXI_READ";
        traffic_data[739].size_bytes = 64;
        traffic_data[740].timestamp = 486;
        traffic_data[740].source_node = 0;
        traffic_data[740].dest_node = 2;
        traffic_data[740].packet_type = "AXI_READ";
        traffic_data[740].size_bytes = 64;
        traffic_data[741].timestamp = 486;
        traffic_data[741].source_node = 7;
        traffic_data[741].dest_node = 14;
        traffic_data[741].packet_type = "CHI_WRITE";
        traffic_data[741].size_bytes = 64;
        traffic_data[742].timestamp = 487;
        traffic_data[742].source_node = 5;
        traffic_data[742].dest_node = 13;
        traffic_data[742].packet_type = "AXI_WRITE";
        traffic_data[742].size_bytes = 64;
        traffic_data[743].timestamp = 487;
        traffic_data[743].source_node = 7;
        traffic_data[743].dest_node = 14;
        traffic_data[743].packet_type = "CHI_WRITE";
        traffic_data[743].size_bytes = 64;
        traffic_data[744].timestamp = 489;
        traffic_data[744].source_node = 6;
        traffic_data[744].dest_node = 10;
        traffic_data[744].packet_type = "CHI_READ";
        traffic_data[744].size_bytes = 64;
        traffic_data[745].timestamp = 489;
        traffic_data[745].source_node = 7;
        traffic_data[745].dest_node = 4;
        traffic_data[745].packet_type = "AXI_WRITE";
        traffic_data[745].size_bytes = 64;
        traffic_data[746].timestamp = 489;
        traffic_data[746].source_node = 9;
        traffic_data[746].dest_node = 10;
        traffic_data[746].packet_type = "AXI_READ";
        traffic_data[746].size_bytes = 64;
        traffic_data[747].timestamp = 489;
        traffic_data[747].source_node = 14;
        traffic_data[747].dest_node = 4;
        traffic_data[747].packet_type = "AXI_READ";
        traffic_data[747].size_bytes = 64;
        traffic_data[748].timestamp = 490;
        traffic_data[748].source_node = 3;
        traffic_data[748].dest_node = 6;
        traffic_data[748].packet_type = "AXI_READ";
        traffic_data[748].size_bytes = 64;
        traffic_data[749].timestamp = 490;
        traffic_data[749].source_node = 5;
        traffic_data[749].dest_node = 6;
        traffic_data[749].packet_type = "CHI_READ";
        traffic_data[749].size_bytes = 64;
        traffic_data[750].timestamp = 491;
        traffic_data[750].source_node = 2;
        traffic_data[750].dest_node = 13;
        traffic_data[750].packet_type = "CHI_WRITE";
        traffic_data[750].size_bytes = 64;
        traffic_data[751].timestamp = 491;
        traffic_data[751].source_node = 5;
        traffic_data[751].dest_node = 2;
        traffic_data[751].packet_type = "AXI_WRITE";
        traffic_data[751].size_bytes = 64;
        traffic_data[752].timestamp = 491;
        traffic_data[752].source_node = 7;
        traffic_data[752].dest_node = 11;
        traffic_data[752].packet_type = "AXI_READ";
        traffic_data[752].size_bytes = 64;
        traffic_data[753].timestamp = 492;
        traffic_data[753].source_node = 9;
        traffic_data[753].dest_node = 12;
        traffic_data[753].packet_type = "CHI_WRITE";
        traffic_data[753].size_bytes = 64;
        traffic_data[754].timestamp = 493;
        traffic_data[754].source_node = 0;
        traffic_data[754].dest_node = 1;
        traffic_data[754].packet_type = "AXI_WRITE";
        traffic_data[754].size_bytes = 64;
        traffic_data[755].timestamp = 493;
        traffic_data[755].source_node = 10;
        traffic_data[755].dest_node = 9;
        traffic_data[755].packet_type = "CHI_READ";
        traffic_data[755].size_bytes = 64;
        traffic_data[756].timestamp = 493;
        traffic_data[756].source_node = 12;
        traffic_data[756].dest_node = 11;
        traffic_data[756].packet_type = "CHI_WRITE";
        traffic_data[756].size_bytes = 64;
        traffic_data[757].timestamp = 494;
        traffic_data[757].source_node = 5;
        traffic_data[757].dest_node = 14;
        traffic_data[757].packet_type = "CHI_READ";
        traffic_data[757].size_bytes = 64;
        traffic_data[758].timestamp = 495;
        traffic_data[758].source_node = 8;
        traffic_data[758].dest_node = 14;
        traffic_data[758].packet_type = "AXI_READ";
        traffic_data[758].size_bytes = 64;
        traffic_data[759].timestamp = 495;
        traffic_data[759].source_node = 12;
        traffic_data[759].dest_node = 6;
        traffic_data[759].packet_type = "CHI_WRITE";
        traffic_data[759].size_bytes = 64;
        traffic_data[760].timestamp = 496;
        traffic_data[760].source_node = 9;
        traffic_data[760].dest_node = 5;
        traffic_data[760].packet_type = "CHI_WRITE";
        traffic_data[760].size_bytes = 64;
        traffic_data[761].timestamp = 497;
        traffic_data[761].source_node = 5;
        traffic_data[761].dest_node = 13;
        traffic_data[761].packet_type = "CHI_READ";
        traffic_data[761].size_bytes = 64;
        traffic_data[762].timestamp = 497;
        traffic_data[762].source_node = 10;
        traffic_data[762].dest_node = 13;
        traffic_data[762].packet_type = "CHI_WRITE";
        traffic_data[762].size_bytes = 64;
        traffic_data[763].timestamp = 497;
        traffic_data[763].source_node = 13;
        traffic_data[763].dest_node = 1;
        traffic_data[763].packet_type = "CHI_READ";
        traffic_data[763].size_bytes = 64;
        traffic_data[764].timestamp = 498;
        traffic_data[764].source_node = 6;
        traffic_data[764].dest_node = 15;
        traffic_data[764].packet_type = "CHI_WRITE";
        traffic_data[764].size_bytes = 64;
        traffic_data[765].timestamp = 499;
        traffic_data[765].source_node = 3;
        traffic_data[765].dest_node = 13;
        traffic_data[765].packet_type = "AXI_WRITE";
        traffic_data[765].size_bytes = 64;
        traffic_data[766].timestamp = 499;
        traffic_data[766].source_node = 4;
        traffic_data[766].dest_node = 11;
        traffic_data[766].packet_type = "AXI_WRITE";
        traffic_data[766].size_bytes = 64;
        traffic_data[767].timestamp = 500;
        traffic_data[767].source_node = 3;
        traffic_data[767].dest_node = 8;
        traffic_data[767].packet_type = "AXI_WRITE";
        traffic_data[767].size_bytes = 64;
        traffic_data[768].timestamp = 500;
        traffic_data[768].source_node = 7;
        traffic_data[768].dest_node = 12;
        traffic_data[768].packet_type = "AXI_WRITE";
        traffic_data[768].size_bytes = 64;
        traffic_data[769].timestamp = 501;
        traffic_data[769].source_node = 0;
        traffic_data[769].dest_node = 14;
        traffic_data[769].packet_type = "CHI_READ";
        traffic_data[769].size_bytes = 64;
        traffic_data[770].timestamp = 501;
        traffic_data[770].source_node = 1;
        traffic_data[770].dest_node = 15;
        traffic_data[770].packet_type = "CHI_READ";
        traffic_data[770].size_bytes = 64;
        traffic_data[771].timestamp = 503;
        traffic_data[771].source_node = 3;
        traffic_data[771].dest_node = 8;
        traffic_data[771].packet_type = "AXI_READ";
        traffic_data[771].size_bytes = 64;
        traffic_data[772].timestamp = 504;
        traffic_data[772].source_node = 12;
        traffic_data[772].dest_node = 15;
        traffic_data[772].packet_type = "CHI_WRITE";
        traffic_data[772].size_bytes = 64;
        traffic_data[773].timestamp = 504;
        traffic_data[773].source_node = 13;
        traffic_data[773].dest_node = 0;
        traffic_data[773].packet_type = "AXI_WRITE";
        traffic_data[773].size_bytes = 64;
        traffic_data[774].timestamp = 505;
        traffic_data[774].source_node = 10;
        traffic_data[774].dest_node = 15;
        traffic_data[774].packet_type = "CHI_WRITE";
        traffic_data[774].size_bytes = 64;
        traffic_data[775].timestamp = 506;
        traffic_data[775].source_node = 2;
        traffic_data[775].dest_node = 13;
        traffic_data[775].packet_type = "AXI_WRITE";
        traffic_data[775].size_bytes = 64;
        traffic_data[776].timestamp = 506;
        traffic_data[776].source_node = 12;
        traffic_data[776].dest_node = 6;
        traffic_data[776].packet_type = "AXI_READ";
        traffic_data[776].size_bytes = 64;
        traffic_data[777].timestamp = 506;
        traffic_data[777].source_node = 15;
        traffic_data[777].dest_node = 11;
        traffic_data[777].packet_type = "AXI_READ";
        traffic_data[777].size_bytes = 64;
        traffic_data[778].timestamp = 507;
        traffic_data[778].source_node = 1;
        traffic_data[778].dest_node = 12;
        traffic_data[778].packet_type = "AXI_WRITE";
        traffic_data[778].size_bytes = 64;
        traffic_data[779].timestamp = 507;
        traffic_data[779].source_node = 14;
        traffic_data[779].dest_node = 1;
        traffic_data[779].packet_type = "AXI_WRITE";
        traffic_data[779].size_bytes = 64;
        traffic_data[780].timestamp = 508;
        traffic_data[780].source_node = 8;
        traffic_data[780].dest_node = 7;
        traffic_data[780].packet_type = "CHI_READ";
        traffic_data[780].size_bytes = 64;
        traffic_data[781].timestamp = 510;
        traffic_data[781].source_node = 0;
        traffic_data[781].dest_node = 9;
        traffic_data[781].packet_type = "CHI_READ";
        traffic_data[781].size_bytes = 64;
        traffic_data[782].timestamp = 510;
        traffic_data[782].source_node = 3;
        traffic_data[782].dest_node = 0;
        traffic_data[782].packet_type = "AXI_WRITE";
        traffic_data[782].size_bytes = 64;
        traffic_data[783].timestamp = 510;
        traffic_data[783].source_node = 7;
        traffic_data[783].dest_node = 2;
        traffic_data[783].packet_type = "AXI_WRITE";
        traffic_data[783].size_bytes = 64;
        traffic_data[784].timestamp = 510;
        traffic_data[784].source_node = 8;
        traffic_data[784].dest_node = 12;
        traffic_data[784].packet_type = "AXI_WRITE";
        traffic_data[784].size_bytes = 64;
        traffic_data[785].timestamp = 512;
        traffic_data[785].source_node = 9;
        traffic_data[785].dest_node = 2;
        traffic_data[785].packet_type = "AXI_READ";
        traffic_data[785].size_bytes = 64;
        traffic_data[786].timestamp = 513;
        traffic_data[786].source_node = 11;
        traffic_data[786].dest_node = 12;
        traffic_data[786].packet_type = "AXI_READ";
        traffic_data[786].size_bytes = 64;
        traffic_data[787].timestamp = 514;
        traffic_data[787].source_node = 1;
        traffic_data[787].dest_node = 5;
        traffic_data[787].packet_type = "AXI_WRITE";
        traffic_data[787].size_bytes = 64;
        traffic_data[788].timestamp = 514;
        traffic_data[788].source_node = 8;
        traffic_data[788].dest_node = 15;
        traffic_data[788].packet_type = "CHI_WRITE";
        traffic_data[788].size_bytes = 64;
        traffic_data[789].timestamp = 514;
        traffic_data[789].source_node = 13;
        traffic_data[789].dest_node = 7;
        traffic_data[789].packet_type = "CHI_WRITE";
        traffic_data[789].size_bytes = 64;
        traffic_data[790].timestamp = 514;
        traffic_data[790].source_node = 14;
        traffic_data[790].dest_node = 4;
        traffic_data[790].packet_type = "CHI_WRITE";
        traffic_data[790].size_bytes = 64;
        traffic_data[791].timestamp = 515;
        traffic_data[791].source_node = 4;
        traffic_data[791].dest_node = 0;
        traffic_data[791].packet_type = "AXI_READ";
        traffic_data[791].size_bytes = 64;
        traffic_data[792].timestamp = 515;
        traffic_data[792].source_node = 11;
        traffic_data[792].dest_node = 10;
        traffic_data[792].packet_type = "AXI_READ";
        traffic_data[792].size_bytes = 64;
        traffic_data[793].timestamp = 515;
        traffic_data[793].source_node = 12;
        traffic_data[793].dest_node = 1;
        traffic_data[793].packet_type = "CHI_WRITE";
        traffic_data[793].size_bytes = 64;
        traffic_data[794].timestamp = 516;
        traffic_data[794].source_node = 12;
        traffic_data[794].dest_node = 0;
        traffic_data[794].packet_type = "AXI_READ";
        traffic_data[794].size_bytes = 64;
        traffic_data[795].timestamp = 517;
        traffic_data[795].source_node = 2;
        traffic_data[795].dest_node = 12;
        traffic_data[795].packet_type = "CHI_READ";
        traffic_data[795].size_bytes = 64;
        traffic_data[796].timestamp = 517;
        traffic_data[796].source_node = 5;
        traffic_data[796].dest_node = 12;
        traffic_data[796].packet_type = "AXI_READ";
        traffic_data[796].size_bytes = 64;
        traffic_data[797].timestamp = 517;
        traffic_data[797].source_node = 10;
        traffic_data[797].dest_node = 5;
        traffic_data[797].packet_type = "CHI_WRITE";
        traffic_data[797].size_bytes = 64;
        traffic_data[798].timestamp = 519;
        traffic_data[798].source_node = 0;
        traffic_data[798].dest_node = 9;
        traffic_data[798].packet_type = "AXI_WRITE";
        traffic_data[798].size_bytes = 64;
        traffic_data[799].timestamp = 519;
        traffic_data[799].source_node = 4;
        traffic_data[799].dest_node = 8;
        traffic_data[799].packet_type = "AXI_READ";
        traffic_data[799].size_bytes = 64;
        traffic_data[800].timestamp = 520;
        traffic_data[800].source_node = 11;
        traffic_data[800].dest_node = 6;
        traffic_data[800].packet_type = "AXI_WRITE";
        traffic_data[800].size_bytes = 64;
        traffic_data[801].timestamp = 521;
        traffic_data[801].source_node = 3;
        traffic_data[801].dest_node = 8;
        traffic_data[801].packet_type = "AXI_WRITE";
        traffic_data[801].size_bytes = 64;
        traffic_data[802].timestamp = 522;
        traffic_data[802].source_node = 1;
        traffic_data[802].dest_node = 7;
        traffic_data[802].packet_type = "CHI_WRITE";
        traffic_data[802].size_bytes = 64;
        traffic_data[803].timestamp = 522;
        traffic_data[803].source_node = 9;
        traffic_data[803].dest_node = 3;
        traffic_data[803].packet_type = "AXI_READ";
        traffic_data[803].size_bytes = 64;
        traffic_data[804].timestamp = 522;
        traffic_data[804].source_node = 11;
        traffic_data[804].dest_node = 0;
        traffic_data[804].packet_type = "CHI_READ";
        traffic_data[804].size_bytes = 64;
        traffic_data[805].timestamp = 523;
        traffic_data[805].source_node = 12;
        traffic_data[805].dest_node = 2;
        traffic_data[805].packet_type = "CHI_WRITE";
        traffic_data[805].size_bytes = 64;
        traffic_data[806].timestamp = 524;
        traffic_data[806].source_node = 8;
        traffic_data[806].dest_node = 4;
        traffic_data[806].packet_type = "AXI_READ";
        traffic_data[806].size_bytes = 64;
        traffic_data[807].timestamp = 524;
        traffic_data[807].source_node = 11;
        traffic_data[807].dest_node = 5;
        traffic_data[807].packet_type = "CHI_WRITE";
        traffic_data[807].size_bytes = 64;
        traffic_data[808].timestamp = 525;
        traffic_data[808].source_node = 7;
        traffic_data[808].dest_node = 4;
        traffic_data[808].packet_type = "CHI_READ";
        traffic_data[808].size_bytes = 64;
        traffic_data[809].timestamp = 525;
        traffic_data[809].source_node = 14;
        traffic_data[809].dest_node = 5;
        traffic_data[809].packet_type = "CHI_READ";
        traffic_data[809].size_bytes = 64;
        traffic_data[810].timestamp = 526;
        traffic_data[810].source_node = 8;
        traffic_data[810].dest_node = 6;
        traffic_data[810].packet_type = "AXI_WRITE";
        traffic_data[810].size_bytes = 64;
        traffic_data[811].timestamp = 528;
        traffic_data[811].source_node = 2;
        traffic_data[811].dest_node = 9;
        traffic_data[811].packet_type = "CHI_READ";
        traffic_data[811].size_bytes = 64;
        traffic_data[812].timestamp = 528;
        traffic_data[812].source_node = 10;
        traffic_data[812].dest_node = 15;
        traffic_data[812].packet_type = "AXI_WRITE";
        traffic_data[812].size_bytes = 64;
        traffic_data[813].timestamp = 529;
        traffic_data[813].source_node = 3;
        traffic_data[813].dest_node = 0;
        traffic_data[813].packet_type = "AXI_WRITE";
        traffic_data[813].size_bytes = 64;
        traffic_data[814].timestamp = 529;
        traffic_data[814].source_node = 6;
        traffic_data[814].dest_node = 4;
        traffic_data[814].packet_type = "AXI_READ";
        traffic_data[814].size_bytes = 64;
        traffic_data[815].timestamp = 529;
        traffic_data[815].source_node = 9;
        traffic_data[815].dest_node = 4;
        traffic_data[815].packet_type = "AXI_WRITE";
        traffic_data[815].size_bytes = 64;
        traffic_data[816].timestamp = 530;
        traffic_data[816].source_node = 0;
        traffic_data[816].dest_node = 5;
        traffic_data[816].packet_type = "AXI_WRITE";
        traffic_data[816].size_bytes = 64;
        traffic_data[817].timestamp = 530;
        traffic_data[817].source_node = 4;
        traffic_data[817].dest_node = 3;
        traffic_data[817].packet_type = "AXI_READ";
        traffic_data[817].size_bytes = 64;
        traffic_data[818].timestamp = 530;
        traffic_data[818].source_node = 11;
        traffic_data[818].dest_node = 4;
        traffic_data[818].packet_type = "CHI_READ";
        traffic_data[818].size_bytes = 64;
        traffic_data[819].timestamp = 531;
        traffic_data[819].source_node = 13;
        traffic_data[819].dest_node = 8;
        traffic_data[819].packet_type = "CHI_WRITE";
        traffic_data[819].size_bytes = 64;
        traffic_data[820].timestamp = 532;
        traffic_data[820].source_node = 7;
        traffic_data[820].dest_node = 13;
        traffic_data[820].packet_type = "CHI_WRITE";
        traffic_data[820].size_bytes = 64;
        traffic_data[821].timestamp = 532;
        traffic_data[821].source_node = 8;
        traffic_data[821].dest_node = 2;
        traffic_data[821].packet_type = "CHI_READ";
        traffic_data[821].size_bytes = 64;
        traffic_data[822].timestamp = 532;
        traffic_data[822].source_node = 15;
        traffic_data[822].dest_node = 13;
        traffic_data[822].packet_type = "CHI_WRITE";
        traffic_data[822].size_bytes = 64;
        traffic_data[823].timestamp = 533;
        traffic_data[823].source_node = 6;
        traffic_data[823].dest_node = 4;
        traffic_data[823].packet_type = "AXI_READ";
        traffic_data[823].size_bytes = 64;
        traffic_data[824].timestamp = 533;
        traffic_data[824].source_node = 8;
        traffic_data[824].dest_node = 4;
        traffic_data[824].packet_type = "CHI_WRITE";
        traffic_data[824].size_bytes = 64;
        traffic_data[825].timestamp = 534;
        traffic_data[825].source_node = 13;
        traffic_data[825].dest_node = 2;
        traffic_data[825].packet_type = "AXI_READ";
        traffic_data[825].size_bytes = 64;
        traffic_data[826].timestamp = 535;
        traffic_data[826].source_node = 1;
        traffic_data[826].dest_node = 9;
        traffic_data[826].packet_type = "CHI_WRITE";
        traffic_data[826].size_bytes = 64;
        traffic_data[827].timestamp = 535;
        traffic_data[827].source_node = 15;
        traffic_data[827].dest_node = 2;
        traffic_data[827].packet_type = "AXI_WRITE";
        traffic_data[827].size_bytes = 64;
        traffic_data[828].timestamp = 536;
        traffic_data[828].source_node = 14;
        traffic_data[828].dest_node = 7;
        traffic_data[828].packet_type = "AXI_READ";
        traffic_data[828].size_bytes = 64;
        traffic_data[829].timestamp = 537;
        traffic_data[829].source_node = 0;
        traffic_data[829].dest_node = 5;
        traffic_data[829].packet_type = "AXI_READ";
        traffic_data[829].size_bytes = 64;
        traffic_data[830].timestamp = 537;
        traffic_data[830].source_node = 4;
        traffic_data[830].dest_node = 15;
        traffic_data[830].packet_type = "CHI_READ";
        traffic_data[830].size_bytes = 64;
        traffic_data[831].timestamp = 538;
        traffic_data[831].source_node = 0;
        traffic_data[831].dest_node = 11;
        traffic_data[831].packet_type = "AXI_WRITE";
        traffic_data[831].size_bytes = 64;
        traffic_data[832].timestamp = 539;
        traffic_data[832].source_node = 9;
        traffic_data[832].dest_node = 14;
        traffic_data[832].packet_type = "AXI_WRITE";
        traffic_data[832].size_bytes = 64;
        traffic_data[833].timestamp = 540;
        traffic_data[833].source_node = 9;
        traffic_data[833].dest_node = 4;
        traffic_data[833].packet_type = "AXI_READ";
        traffic_data[833].size_bytes = 64;
        traffic_data[834].timestamp = 540;
        traffic_data[834].source_node = 10;
        traffic_data[834].dest_node = 12;
        traffic_data[834].packet_type = "AXI_READ";
        traffic_data[834].size_bytes = 64;
        traffic_data[835].timestamp = 540;
        traffic_data[835].source_node = 14;
        traffic_data[835].dest_node = 2;
        traffic_data[835].packet_type = "CHI_READ";
        traffic_data[835].size_bytes = 64;
        traffic_data[836].timestamp = 541;
        traffic_data[836].source_node = 12;
        traffic_data[836].dest_node = 0;
        traffic_data[836].packet_type = "AXI_READ";
        traffic_data[836].size_bytes = 64;
        traffic_data[837].timestamp = 542;
        traffic_data[837].source_node = 3;
        traffic_data[837].dest_node = 2;
        traffic_data[837].packet_type = "CHI_WRITE";
        traffic_data[837].size_bytes = 64;
        traffic_data[838].timestamp = 543;
        traffic_data[838].source_node = 4;
        traffic_data[838].dest_node = 9;
        traffic_data[838].packet_type = "CHI_READ";
        traffic_data[838].size_bytes = 64;
        traffic_data[839].timestamp = 543;
        traffic_data[839].source_node = 5;
        traffic_data[839].dest_node = 14;
        traffic_data[839].packet_type = "CHI_READ";
        traffic_data[839].size_bytes = 64;
        traffic_data[840].timestamp = 543;
        traffic_data[840].source_node = 9;
        traffic_data[840].dest_node = 14;
        traffic_data[840].packet_type = "AXI_WRITE";
        traffic_data[840].size_bytes = 64;
        traffic_data[841].timestamp = 543;
        traffic_data[841].source_node = 11;
        traffic_data[841].dest_node = 9;
        traffic_data[841].packet_type = "AXI_WRITE";
        traffic_data[841].size_bytes = 64;
        traffic_data[842].timestamp = 544;
        traffic_data[842].source_node = 0;
        traffic_data[842].dest_node = 12;
        traffic_data[842].packet_type = "AXI_READ";
        traffic_data[842].size_bytes = 64;
        traffic_data[843].timestamp = 544;
        traffic_data[843].source_node = 5;
        traffic_data[843].dest_node = 7;
        traffic_data[843].packet_type = "CHI_READ";
        traffic_data[843].size_bytes = 64;
        traffic_data[844].timestamp = 544;
        traffic_data[844].source_node = 8;
        traffic_data[844].dest_node = 3;
        traffic_data[844].packet_type = "CHI_READ";
        traffic_data[844].size_bytes = 64;
        traffic_data[845].timestamp = 544;
        traffic_data[845].source_node = 13;
        traffic_data[845].dest_node = 9;
        traffic_data[845].packet_type = "AXI_READ";
        traffic_data[845].size_bytes = 64;
        traffic_data[846].timestamp = 544;
        traffic_data[846].source_node = 15;
        traffic_data[846].dest_node = 6;
        traffic_data[846].packet_type = "AXI_READ";
        traffic_data[846].size_bytes = 64;
        traffic_data[847].timestamp = 545;
        traffic_data[847].source_node = 13;
        traffic_data[847].dest_node = 12;
        traffic_data[847].packet_type = "AXI_WRITE";
        traffic_data[847].size_bytes = 64;
        traffic_data[848].timestamp = 546;
        traffic_data[848].source_node = 3;
        traffic_data[848].dest_node = 13;
        traffic_data[848].packet_type = "CHI_WRITE";
        traffic_data[848].size_bytes = 64;
        traffic_data[849].timestamp = 546;
        traffic_data[849].source_node = 14;
        traffic_data[849].dest_node = 3;
        traffic_data[849].packet_type = "AXI_READ";
        traffic_data[849].size_bytes = 64;
        traffic_data[850].timestamp = 547;
        traffic_data[850].source_node = 6;
        traffic_data[850].dest_node = 12;
        traffic_data[850].packet_type = "AXI_WRITE";
        traffic_data[850].size_bytes = 64;
        traffic_data[851].timestamp = 547;
        traffic_data[851].source_node = 8;
        traffic_data[851].dest_node = 2;
        traffic_data[851].packet_type = "CHI_WRITE";
        traffic_data[851].size_bytes = 64;
        traffic_data[852].timestamp = 547;
        traffic_data[852].source_node = 10;
        traffic_data[852].dest_node = 5;
        traffic_data[852].packet_type = "AXI_WRITE";
        traffic_data[852].size_bytes = 64;
        traffic_data[853].timestamp = 548;
        traffic_data[853].source_node = 0;
        traffic_data[853].dest_node = 9;
        traffic_data[853].packet_type = "AXI_WRITE";
        traffic_data[853].size_bytes = 64;
        traffic_data[854].timestamp = 548;
        traffic_data[854].source_node = 15;
        traffic_data[854].dest_node = 14;
        traffic_data[854].packet_type = "CHI_WRITE";
        traffic_data[854].size_bytes = 64;
        traffic_data[855].timestamp = 550;
        traffic_data[855].source_node = 2;
        traffic_data[855].dest_node = 5;
        traffic_data[855].packet_type = "CHI_WRITE";
        traffic_data[855].size_bytes = 64;
        traffic_data[856].timestamp = 550;
        traffic_data[856].source_node = 5;
        traffic_data[856].dest_node = 14;
        traffic_data[856].packet_type = "CHI_WRITE";
        traffic_data[856].size_bytes = 64;
        traffic_data[857].timestamp = 550;
        traffic_data[857].source_node = 9;
        traffic_data[857].dest_node = 3;
        traffic_data[857].packet_type = "CHI_WRITE";
        traffic_data[857].size_bytes = 64;
        traffic_data[858].timestamp = 550;
        traffic_data[858].source_node = 12;
        traffic_data[858].dest_node = 4;
        traffic_data[858].packet_type = "AXI_READ";
        traffic_data[858].size_bytes = 64;
        traffic_data[859].timestamp = 550;
        traffic_data[859].source_node = 15;
        traffic_data[859].dest_node = 9;
        traffic_data[859].packet_type = "CHI_READ";
        traffic_data[859].size_bytes = 64;
        traffic_data[860].timestamp = 551;
        traffic_data[860].source_node = 11;
        traffic_data[860].dest_node = 1;
        traffic_data[860].packet_type = "CHI_WRITE";
        traffic_data[860].size_bytes = 64;
        traffic_data[861].timestamp = 553;
        traffic_data[861].source_node = 1;
        traffic_data[861].dest_node = 5;
        traffic_data[861].packet_type = "CHI_READ";
        traffic_data[861].size_bytes = 64;
        traffic_data[862].timestamp = 553;
        traffic_data[862].source_node = 6;
        traffic_data[862].dest_node = 4;
        traffic_data[862].packet_type = "CHI_READ";
        traffic_data[862].size_bytes = 64;
        traffic_data[863].timestamp = 553;
        traffic_data[863].source_node = 10;
        traffic_data[863].dest_node = 0;
        traffic_data[863].packet_type = "CHI_WRITE";
        traffic_data[863].size_bytes = 64;
        traffic_data[864].timestamp = 553;
        traffic_data[864].source_node = 11;
        traffic_data[864].dest_node = 5;
        traffic_data[864].packet_type = "CHI_WRITE";
        traffic_data[864].size_bytes = 64;
        traffic_data[865].timestamp = 554;
        traffic_data[865].source_node = 0;
        traffic_data[865].dest_node = 15;
        traffic_data[865].packet_type = "CHI_READ";
        traffic_data[865].size_bytes = 64;
        traffic_data[866].timestamp = 555;
        traffic_data[866].source_node = 6;
        traffic_data[866].dest_node = 14;
        traffic_data[866].packet_type = "CHI_READ";
        traffic_data[866].size_bytes = 64;
        traffic_data[867].timestamp = 555;
        traffic_data[867].source_node = 8;
        traffic_data[867].dest_node = 3;
        traffic_data[867].packet_type = "CHI_READ";
        traffic_data[867].size_bytes = 64;
        traffic_data[868].timestamp = 555;
        traffic_data[868].source_node = 12;
        traffic_data[868].dest_node = 3;
        traffic_data[868].packet_type = "CHI_READ";
        traffic_data[868].size_bytes = 64;
        traffic_data[869].timestamp = 556;
        traffic_data[869].source_node = 0;
        traffic_data[869].dest_node = 7;
        traffic_data[869].packet_type = "CHI_READ";
        traffic_data[869].size_bytes = 64;
        traffic_data[870].timestamp = 556;
        traffic_data[870].source_node = 11;
        traffic_data[870].dest_node = 15;
        traffic_data[870].packet_type = "AXI_WRITE";
        traffic_data[870].size_bytes = 64;
        traffic_data[871].timestamp = 556;
        traffic_data[871].source_node = 13;
        traffic_data[871].dest_node = 9;
        traffic_data[871].packet_type = "AXI_WRITE";
        traffic_data[871].size_bytes = 64;
        traffic_data[872].timestamp = 557;
        traffic_data[872].source_node = 6;
        traffic_data[872].dest_node = 12;
        traffic_data[872].packet_type = "AXI_WRITE";
        traffic_data[872].size_bytes = 64;
        traffic_data[873].timestamp = 557;
        traffic_data[873].source_node = 9;
        traffic_data[873].dest_node = 1;
        traffic_data[873].packet_type = "AXI_WRITE";
        traffic_data[873].size_bytes = 64;
        traffic_data[874].timestamp = 559;
        traffic_data[874].source_node = 3;
        traffic_data[874].dest_node = 9;
        traffic_data[874].packet_type = "AXI_READ";
        traffic_data[874].size_bytes = 64;
        traffic_data[875].timestamp = 560;
        traffic_data[875].source_node = 4;
        traffic_data[875].dest_node = 7;
        traffic_data[875].packet_type = "AXI_WRITE";
        traffic_data[875].size_bytes = 64;
        traffic_data[876].timestamp = 560;
        traffic_data[876].source_node = 10;
        traffic_data[876].dest_node = 1;
        traffic_data[876].packet_type = "CHI_WRITE";
        traffic_data[876].size_bytes = 64;
        traffic_data[877].timestamp = 561;
        traffic_data[877].source_node = 0;
        traffic_data[877].dest_node = 7;
        traffic_data[877].packet_type = "AXI_READ";
        traffic_data[877].size_bytes = 64;
        traffic_data[878].timestamp = 562;
        traffic_data[878].source_node = 1;
        traffic_data[878].dest_node = 12;
        traffic_data[878].packet_type = "CHI_READ";
        traffic_data[878].size_bytes = 64;
        traffic_data[879].timestamp = 562;
        traffic_data[879].source_node = 15;
        traffic_data[879].dest_node = 9;
        traffic_data[879].packet_type = "CHI_READ";
        traffic_data[879].size_bytes = 64;
        traffic_data[880].timestamp = 563;
        traffic_data[880].source_node = 9;
        traffic_data[880].dest_node = 8;
        traffic_data[880].packet_type = "CHI_WRITE";
        traffic_data[880].size_bytes = 64;
        traffic_data[881].timestamp = 563;
        traffic_data[881].source_node = 14;
        traffic_data[881].dest_node = 11;
        traffic_data[881].packet_type = "AXI_WRITE";
        traffic_data[881].size_bytes = 64;
        traffic_data[882].timestamp = 564;
        traffic_data[882].source_node = 15;
        traffic_data[882].dest_node = 8;
        traffic_data[882].packet_type = "AXI_WRITE";
        traffic_data[882].size_bytes = 64;
        traffic_data[883].timestamp = 565;
        traffic_data[883].source_node = 0;
        traffic_data[883].dest_node = 15;
        traffic_data[883].packet_type = "AXI_READ";
        traffic_data[883].size_bytes = 64;
        traffic_data[884].timestamp = 565;
        traffic_data[884].source_node = 4;
        traffic_data[884].dest_node = 14;
        traffic_data[884].packet_type = "AXI_READ";
        traffic_data[884].size_bytes = 64;
        traffic_data[885].timestamp = 566;
        traffic_data[885].source_node = 2;
        traffic_data[885].dest_node = 3;
        traffic_data[885].packet_type = "CHI_READ";
        traffic_data[885].size_bytes = 64;
        traffic_data[886].timestamp = 566;
        traffic_data[886].source_node = 6;
        traffic_data[886].dest_node = 13;
        traffic_data[886].packet_type = "AXI_WRITE";
        traffic_data[886].size_bytes = 64;
        traffic_data[887].timestamp = 567;
        traffic_data[887].source_node = 8;
        traffic_data[887].dest_node = 11;
        traffic_data[887].packet_type = "AXI_READ";
        traffic_data[887].size_bytes = 64;
        traffic_data[888].timestamp = 568;
        traffic_data[888].source_node = 4;
        traffic_data[888].dest_node = 9;
        traffic_data[888].packet_type = "AXI_WRITE";
        traffic_data[888].size_bytes = 64;
        traffic_data[889].timestamp = 568;
        traffic_data[889].source_node = 5;
        traffic_data[889].dest_node = 1;
        traffic_data[889].packet_type = "CHI_WRITE";
        traffic_data[889].size_bytes = 64;
        traffic_data[890].timestamp = 569;
        traffic_data[890].source_node = 9;
        traffic_data[890].dest_node = 1;
        traffic_data[890].packet_type = "CHI_READ";
        traffic_data[890].size_bytes = 64;
        traffic_data[891].timestamp = 570;
        traffic_data[891].source_node = 9;
        traffic_data[891].dest_node = 4;
        traffic_data[891].packet_type = "AXI_WRITE";
        traffic_data[891].size_bytes = 64;
        traffic_data[892].timestamp = 570;
        traffic_data[892].source_node = 12;
        traffic_data[892].dest_node = 13;
        traffic_data[892].packet_type = "CHI_READ";
        traffic_data[892].size_bytes = 64;
        traffic_data[893].timestamp = 572;
        traffic_data[893].source_node = 1;
        traffic_data[893].dest_node = 12;
        traffic_data[893].packet_type = "AXI_READ";
        traffic_data[893].size_bytes = 64;
        traffic_data[894].timestamp = 572;
        traffic_data[894].source_node = 3;
        traffic_data[894].dest_node = 12;
        traffic_data[894].packet_type = "CHI_READ";
        traffic_data[894].size_bytes = 64;
        traffic_data[895].timestamp = 573;
        traffic_data[895].source_node = 5;
        traffic_data[895].dest_node = 0;
        traffic_data[895].packet_type = "AXI_READ";
        traffic_data[895].size_bytes = 64;
        traffic_data[896].timestamp = 573;
        traffic_data[896].source_node = 8;
        traffic_data[896].dest_node = 4;
        traffic_data[896].packet_type = "CHI_READ";
        traffic_data[896].size_bytes = 64;
        traffic_data[897].timestamp = 573;
        traffic_data[897].source_node = 9;
        traffic_data[897].dest_node = 11;
        traffic_data[897].packet_type = "AXI_WRITE";
        traffic_data[897].size_bytes = 64;
        traffic_data[898].timestamp = 573;
        traffic_data[898].source_node = 10;
        traffic_data[898].dest_node = 12;
        traffic_data[898].packet_type = "AXI_READ";
        traffic_data[898].size_bytes = 64;
        traffic_data[899].timestamp = 574;
        traffic_data[899].source_node = 1;
        traffic_data[899].dest_node = 9;
        traffic_data[899].packet_type = "CHI_WRITE";
        traffic_data[899].size_bytes = 64;
        traffic_data[900].timestamp = 574;
        traffic_data[900].source_node = 2;
        traffic_data[900].dest_node = 12;
        traffic_data[900].packet_type = "AXI_WRITE";
        traffic_data[900].size_bytes = 64;
        traffic_data[901].timestamp = 574;
        traffic_data[901].source_node = 3;
        traffic_data[901].dest_node = 10;
        traffic_data[901].packet_type = "CHI_WRITE";
        traffic_data[901].size_bytes = 64;
        traffic_data[902].timestamp = 574;
        traffic_data[902].source_node = 9;
        traffic_data[902].dest_node = 4;
        traffic_data[902].packet_type = "CHI_WRITE";
        traffic_data[902].size_bytes = 64;
        traffic_data[903].timestamp = 574;
        traffic_data[903].source_node = 15;
        traffic_data[903].dest_node = 6;
        traffic_data[903].packet_type = "CHI_READ";
        traffic_data[903].size_bytes = 64;
        traffic_data[904].timestamp = 575;
        traffic_data[904].source_node = 4;
        traffic_data[904].dest_node = 8;
        traffic_data[904].packet_type = "CHI_WRITE";
        traffic_data[904].size_bytes = 64;
        traffic_data[905].timestamp = 575;
        traffic_data[905].source_node = 10;
        traffic_data[905].dest_node = 13;
        traffic_data[905].packet_type = "AXI_WRITE";
        traffic_data[905].size_bytes = 64;
        traffic_data[906].timestamp = 576;
        traffic_data[906].source_node = 1;
        traffic_data[906].dest_node = 9;
        traffic_data[906].packet_type = "AXI_WRITE";
        traffic_data[906].size_bytes = 64;
        traffic_data[907].timestamp = 576;
        traffic_data[907].source_node = 5;
        traffic_data[907].dest_node = 7;
        traffic_data[907].packet_type = "CHI_WRITE";
        traffic_data[907].size_bytes = 64;
        traffic_data[908].timestamp = 576;
        traffic_data[908].source_node = 9;
        traffic_data[908].dest_node = 7;
        traffic_data[908].packet_type = "CHI_READ";
        traffic_data[908].size_bytes = 64;
        traffic_data[909].timestamp = 576;
        traffic_data[909].source_node = 13;
        traffic_data[909].dest_node = 11;
        traffic_data[909].packet_type = "CHI_WRITE";
        traffic_data[909].size_bytes = 64;
        traffic_data[910].timestamp = 577;
        traffic_data[910].source_node = 13;
        traffic_data[910].dest_node = 2;
        traffic_data[910].packet_type = "AXI_READ";
        traffic_data[910].size_bytes = 64;
        traffic_data[911].timestamp = 578;
        traffic_data[911].source_node = 3;
        traffic_data[911].dest_node = 7;
        traffic_data[911].packet_type = "CHI_WRITE";
        traffic_data[911].size_bytes = 64;
        traffic_data[912].timestamp = 580;
        traffic_data[912].source_node = 2;
        traffic_data[912].dest_node = 7;
        traffic_data[912].packet_type = "AXI_WRITE";
        traffic_data[912].size_bytes = 64;
        traffic_data[913].timestamp = 580;
        traffic_data[913].source_node = 4;
        traffic_data[913].dest_node = 0;
        traffic_data[913].packet_type = "CHI_READ";
        traffic_data[913].size_bytes = 64;
        traffic_data[914].timestamp = 580;
        traffic_data[914].source_node = 7;
        traffic_data[914].dest_node = 8;
        traffic_data[914].packet_type = "CHI_READ";
        traffic_data[914].size_bytes = 64;
        traffic_data[915].timestamp = 580;
        traffic_data[915].source_node = 8;
        traffic_data[915].dest_node = 10;
        traffic_data[915].packet_type = "CHI_WRITE";
        traffic_data[915].size_bytes = 64;
        traffic_data[916].timestamp = 580;
        traffic_data[916].source_node = 10;
        traffic_data[916].dest_node = 11;
        traffic_data[916].packet_type = "AXI_WRITE";
        traffic_data[916].size_bytes = 64;
        traffic_data[917].timestamp = 580;
        traffic_data[917].source_node = 12;
        traffic_data[917].dest_node = 3;
        traffic_data[917].packet_type = "CHI_READ";
        traffic_data[917].size_bytes = 64;
        traffic_data[918].timestamp = 582;
        traffic_data[918].source_node = 8;
        traffic_data[918].dest_node = 3;
        traffic_data[918].packet_type = "AXI_WRITE";
        traffic_data[918].size_bytes = 64;
        traffic_data[919].timestamp = 582;
        traffic_data[919].source_node = 9;
        traffic_data[919].dest_node = 13;
        traffic_data[919].packet_type = "AXI_WRITE";
        traffic_data[919].size_bytes = 64;
        traffic_data[920].timestamp = 582;
        traffic_data[920].source_node = 12;
        traffic_data[920].dest_node = 1;
        traffic_data[920].packet_type = "AXI_READ";
        traffic_data[920].size_bytes = 64;
        traffic_data[921].timestamp = 583;
        traffic_data[921].source_node = 10;
        traffic_data[921].dest_node = 9;
        traffic_data[921].packet_type = "AXI_WRITE";
        traffic_data[921].size_bytes = 64;
        traffic_data[922].timestamp = 584;
        traffic_data[922].source_node = 7;
        traffic_data[922].dest_node = 5;
        traffic_data[922].packet_type = "CHI_WRITE";
        traffic_data[922].size_bytes = 64;
        traffic_data[923].timestamp = 585;
        traffic_data[923].source_node = 10;
        traffic_data[923].dest_node = 4;
        traffic_data[923].packet_type = "AXI_READ";
        traffic_data[923].size_bytes = 64;
        traffic_data[924].timestamp = 586;
        traffic_data[924].source_node = 1;
        traffic_data[924].dest_node = 10;
        traffic_data[924].packet_type = "AXI_READ";
        traffic_data[924].size_bytes = 64;
        traffic_data[925].timestamp = 586;
        traffic_data[925].source_node = 11;
        traffic_data[925].dest_node = 0;
        traffic_data[925].packet_type = "AXI_WRITE";
        traffic_data[925].size_bytes = 64;
        traffic_data[926].timestamp = 586;
        traffic_data[926].source_node = 15;
        traffic_data[926].dest_node = 13;
        traffic_data[926].packet_type = "AXI_READ";
        traffic_data[926].size_bytes = 64;
        traffic_data[927].timestamp = 587;
        traffic_data[927].source_node = 0;
        traffic_data[927].dest_node = 11;
        traffic_data[927].packet_type = "AXI_READ";
        traffic_data[927].size_bytes = 64;
        traffic_data[928].timestamp = 587;
        traffic_data[928].source_node = 15;
        traffic_data[928].dest_node = 10;
        traffic_data[928].packet_type = "CHI_WRITE";
        traffic_data[928].size_bytes = 64;
        traffic_data[929].timestamp = 588;
        traffic_data[929].source_node = 2;
        traffic_data[929].dest_node = 4;
        traffic_data[929].packet_type = "AXI_WRITE";
        traffic_data[929].size_bytes = 64;
        traffic_data[930].timestamp = 588;
        traffic_data[930].source_node = 4;
        traffic_data[930].dest_node = 8;
        traffic_data[930].packet_type = "AXI_READ";
        traffic_data[930].size_bytes = 64;
        traffic_data[931].timestamp = 588;
        traffic_data[931].source_node = 11;
        traffic_data[931].dest_node = 4;
        traffic_data[931].packet_type = "CHI_READ";
        traffic_data[931].size_bytes = 64;
        traffic_data[932].timestamp = 588;
        traffic_data[932].source_node = 15;
        traffic_data[932].dest_node = 14;
        traffic_data[932].packet_type = "CHI_WRITE";
        traffic_data[932].size_bytes = 64;
        traffic_data[933].timestamp = 589;
        traffic_data[933].source_node = 0;
        traffic_data[933].dest_node = 15;
        traffic_data[933].packet_type = "AXI_READ";
        traffic_data[933].size_bytes = 64;
        traffic_data[934].timestamp = 589;
        traffic_data[934].source_node = 2;
        traffic_data[934].dest_node = 6;
        traffic_data[934].packet_type = "AXI_READ";
        traffic_data[934].size_bytes = 64;
        traffic_data[935].timestamp = 589;
        traffic_data[935].source_node = 7;
        traffic_data[935].dest_node = 12;
        traffic_data[935].packet_type = "AXI_WRITE";
        traffic_data[935].size_bytes = 64;
        traffic_data[936].timestamp = 590;
        traffic_data[936].source_node = 10;
        traffic_data[936].dest_node = 5;
        traffic_data[936].packet_type = "CHI_READ";
        traffic_data[936].size_bytes = 64;
        traffic_data[937].timestamp = 591;
        traffic_data[937].source_node = 0;
        traffic_data[937].dest_node = 14;
        traffic_data[937].packet_type = "CHI_WRITE";
        traffic_data[937].size_bytes = 64;
        traffic_data[938].timestamp = 594;
        traffic_data[938].source_node = 2;
        traffic_data[938].dest_node = 15;
        traffic_data[938].packet_type = "AXI_WRITE";
        traffic_data[938].size_bytes = 64;
        traffic_data[939].timestamp = 594;
        traffic_data[939].source_node = 10;
        traffic_data[939].dest_node = 8;
        traffic_data[939].packet_type = "AXI_WRITE";
        traffic_data[939].size_bytes = 64;
        traffic_data[940].timestamp = 595;
        traffic_data[940].source_node = 11;
        traffic_data[940].dest_node = 2;
        traffic_data[940].packet_type = "AXI_WRITE";
        traffic_data[940].size_bytes = 64;
        traffic_data[941].timestamp = 595;
        traffic_data[941].source_node = 14;
        traffic_data[941].dest_node = 3;
        traffic_data[941].packet_type = "AXI_WRITE";
        traffic_data[941].size_bytes = 64;
        traffic_data[942].timestamp = 596;
        traffic_data[942].source_node = 4;
        traffic_data[942].dest_node = 2;
        traffic_data[942].packet_type = "CHI_READ";
        traffic_data[942].size_bytes = 64;
        traffic_data[943].timestamp = 596;
        traffic_data[943].source_node = 5;
        traffic_data[943].dest_node = 9;
        traffic_data[943].packet_type = "CHI_WRITE";
        traffic_data[943].size_bytes = 64;
        traffic_data[944].timestamp = 596;
        traffic_data[944].source_node = 12;
        traffic_data[944].dest_node = 2;
        traffic_data[944].packet_type = "CHI_READ";
        traffic_data[944].size_bytes = 64;
        traffic_data[945].timestamp = 597;
        traffic_data[945].source_node = 5;
        traffic_data[945].dest_node = 8;
        traffic_data[945].packet_type = "AXI_READ";
        traffic_data[945].size_bytes = 64;
        traffic_data[946].timestamp = 598;
        traffic_data[946].source_node = 10;
        traffic_data[946].dest_node = 6;
        traffic_data[946].packet_type = "AXI_WRITE";
        traffic_data[946].size_bytes = 64;
        traffic_data[947].timestamp = 598;
        traffic_data[947].source_node = 15;
        traffic_data[947].dest_node = 10;
        traffic_data[947].packet_type = "AXI_READ";
        traffic_data[947].size_bytes = 64;
        traffic_data[948].timestamp = 599;
        traffic_data[948].source_node = 7;
        traffic_data[948].dest_node = 11;
        traffic_data[948].packet_type = "CHI_WRITE";
        traffic_data[948].size_bytes = 64;
        traffic_data[949].timestamp = 599;
        traffic_data[949].source_node = 9;
        traffic_data[949].dest_node = 6;
        traffic_data[949].packet_type = "CHI_READ";
        traffic_data[949].size_bytes = 64;
        traffic_data[950].timestamp = 600;
        traffic_data[950].source_node = 8;
        traffic_data[950].dest_node = 0;
        traffic_data[950].packet_type = "CHI_READ";
        traffic_data[950].size_bytes = 64;
        traffic_data[951].timestamp = 601;
        traffic_data[951].source_node = 1;
        traffic_data[951].dest_node = 14;
        traffic_data[951].packet_type = "CHI_WRITE";
        traffic_data[951].size_bytes = 64;
        traffic_data[952].timestamp = 601;
        traffic_data[952].source_node = 3;
        traffic_data[952].dest_node = 10;
        traffic_data[952].packet_type = "CHI_READ";
        traffic_data[952].size_bytes = 64;
        traffic_data[953].timestamp = 601;
        traffic_data[953].source_node = 11;
        traffic_data[953].dest_node = 5;
        traffic_data[953].packet_type = "CHI_READ";
        traffic_data[953].size_bytes = 64;
        traffic_data[954].timestamp = 601;
        traffic_data[954].source_node = 15;
        traffic_data[954].dest_node = 11;
        traffic_data[954].packet_type = "CHI_WRITE";
        traffic_data[954].size_bytes = 64;
        traffic_data[955].timestamp = 602;
        traffic_data[955].source_node = 1;
        traffic_data[955].dest_node = 2;
        traffic_data[955].packet_type = "AXI_WRITE";
        traffic_data[955].size_bytes = 64;
        traffic_data[956].timestamp = 602;
        traffic_data[956].source_node = 14;
        traffic_data[956].dest_node = 5;
        traffic_data[956].packet_type = "AXI_READ";
        traffic_data[956].size_bytes = 64;
        traffic_data[957].timestamp = 603;
        traffic_data[957].source_node = 5;
        traffic_data[957].dest_node = 15;
        traffic_data[957].packet_type = "CHI_READ";
        traffic_data[957].size_bytes = 64;
        traffic_data[958].timestamp = 603;
        traffic_data[958].source_node = 7;
        traffic_data[958].dest_node = 12;
        traffic_data[958].packet_type = "CHI_READ";
        traffic_data[958].size_bytes = 64;
        traffic_data[959].timestamp = 603;
        traffic_data[959].source_node = 10;
        traffic_data[959].dest_node = 15;
        traffic_data[959].packet_type = "CHI_WRITE";
        traffic_data[959].size_bytes = 64;
        traffic_data[960].timestamp = 604;
        traffic_data[960].source_node = 3;
        traffic_data[960].dest_node = 10;
        traffic_data[960].packet_type = "CHI_WRITE";
        traffic_data[960].size_bytes = 64;
        traffic_data[961].timestamp = 604;
        traffic_data[961].source_node = 10;
        traffic_data[961].dest_node = 6;
        traffic_data[961].packet_type = "AXI_WRITE";
        traffic_data[961].size_bytes = 64;
        traffic_data[962].timestamp = 604;
        traffic_data[962].source_node = 14;
        traffic_data[962].dest_node = 6;
        traffic_data[962].packet_type = "AXI_WRITE";
        traffic_data[962].size_bytes = 64;
        traffic_data[963].timestamp = 605;
        traffic_data[963].source_node = 3;
        traffic_data[963].dest_node = 4;
        traffic_data[963].packet_type = "AXI_READ";
        traffic_data[963].size_bytes = 64;
        traffic_data[964].timestamp = 606;
        traffic_data[964].source_node = 11;
        traffic_data[964].dest_node = 7;
        traffic_data[964].packet_type = "CHI_READ";
        traffic_data[964].size_bytes = 64;
        traffic_data[965].timestamp = 606;
        traffic_data[965].source_node = 12;
        traffic_data[965].dest_node = 11;
        traffic_data[965].packet_type = "CHI_READ";
        traffic_data[965].size_bytes = 64;
        traffic_data[966].timestamp = 609;
        traffic_data[966].source_node = 13;
        traffic_data[966].dest_node = 14;
        traffic_data[966].packet_type = "CHI_READ";
        traffic_data[966].size_bytes = 64;
        traffic_data[967].timestamp = 610;
        traffic_data[967].source_node = 1;
        traffic_data[967].dest_node = 10;
        traffic_data[967].packet_type = "CHI_WRITE";
        traffic_data[967].size_bytes = 64;
        traffic_data[968].timestamp = 611;
        traffic_data[968].source_node = 0;
        traffic_data[968].dest_node = 6;
        traffic_data[968].packet_type = "AXI_READ";
        traffic_data[968].size_bytes = 64;
        traffic_data[969].timestamp = 612;
        traffic_data[969].source_node = 15;
        traffic_data[969].dest_node = 0;
        traffic_data[969].packet_type = "CHI_WRITE";
        traffic_data[969].size_bytes = 64;
        traffic_data[970].timestamp = 613;
        traffic_data[970].source_node = 3;
        traffic_data[970].dest_node = 7;
        traffic_data[970].packet_type = "CHI_READ";
        traffic_data[970].size_bytes = 64;
        traffic_data[971].timestamp = 613;
        traffic_data[971].source_node = 12;
        traffic_data[971].dest_node = 13;
        traffic_data[971].packet_type = "CHI_WRITE";
        traffic_data[971].size_bytes = 64;
        traffic_data[972].timestamp = 613;
        traffic_data[972].source_node = 15;
        traffic_data[972].dest_node = 6;
        traffic_data[972].packet_type = "CHI_WRITE";
        traffic_data[972].size_bytes = 64;
        traffic_data[973].timestamp = 614;
        traffic_data[973].source_node = 13;
        traffic_data[973].dest_node = 10;
        traffic_data[973].packet_type = "AXI_READ";
        traffic_data[973].size_bytes = 64;
        traffic_data[974].timestamp = 615;
        traffic_data[974].source_node = 8;
        traffic_data[974].dest_node = 2;
        traffic_data[974].packet_type = "AXI_WRITE";
        traffic_data[974].size_bytes = 64;
        traffic_data[975].timestamp = 615;
        traffic_data[975].source_node = 10;
        traffic_data[975].dest_node = 15;
        traffic_data[975].packet_type = "CHI_READ";
        traffic_data[975].size_bytes = 64;
        traffic_data[976].timestamp = 616;
        traffic_data[976].source_node = 13;
        traffic_data[976].dest_node = 5;
        traffic_data[976].packet_type = "CHI_WRITE";
        traffic_data[976].size_bytes = 64;
        traffic_data[977].timestamp = 617;
        traffic_data[977].source_node = 13;
        traffic_data[977].dest_node = 3;
        traffic_data[977].packet_type = "CHI_READ";
        traffic_data[977].size_bytes = 64;
        traffic_data[978].timestamp = 618;
        traffic_data[978].source_node = 7;
        traffic_data[978].dest_node = 12;
        traffic_data[978].packet_type = "AXI_WRITE";
        traffic_data[978].size_bytes = 64;
        traffic_data[979].timestamp = 618;
        traffic_data[979].source_node = 10;
        traffic_data[979].dest_node = 11;
        traffic_data[979].packet_type = "AXI_READ";
        traffic_data[979].size_bytes = 64;
        traffic_data[980].timestamp = 619;
        traffic_data[980].source_node = 1;
        traffic_data[980].dest_node = 13;
        traffic_data[980].packet_type = "AXI_READ";
        traffic_data[980].size_bytes = 64;
        traffic_data[981].timestamp = 620;
        traffic_data[981].source_node = 9;
        traffic_data[981].dest_node = 15;
        traffic_data[981].packet_type = "AXI_READ";
        traffic_data[981].size_bytes = 64;
        traffic_data[982].timestamp = 620;
        traffic_data[982].source_node = 14;
        traffic_data[982].dest_node = 3;
        traffic_data[982].packet_type = "AXI_READ";
        traffic_data[982].size_bytes = 64;
        traffic_data[983].timestamp = 621;
        traffic_data[983].source_node = 12;
        traffic_data[983].dest_node = 13;
        traffic_data[983].packet_type = "CHI_WRITE";
        traffic_data[983].size_bytes = 64;
        traffic_data[984].timestamp = 623;
        traffic_data[984].source_node = 1;
        traffic_data[984].dest_node = 7;
        traffic_data[984].packet_type = "CHI_READ";
        traffic_data[984].size_bytes = 64;
        traffic_data[985].timestamp = 623;
        traffic_data[985].source_node = 2;
        traffic_data[985].dest_node = 14;
        traffic_data[985].packet_type = "CHI_WRITE";
        traffic_data[985].size_bytes = 64;
        traffic_data[986].timestamp = 625;
        traffic_data[986].source_node = 9;
        traffic_data[986].dest_node = 6;
        traffic_data[986].packet_type = "AXI_READ";
        traffic_data[986].size_bytes = 64;
        traffic_data[987].timestamp = 625;
        traffic_data[987].source_node = 15;
        traffic_data[987].dest_node = 11;
        traffic_data[987].packet_type = "AXI_WRITE";
        traffic_data[987].size_bytes = 64;
        traffic_data[988].timestamp = 627;
        traffic_data[988].source_node = 3;
        traffic_data[988].dest_node = 11;
        traffic_data[988].packet_type = "CHI_WRITE";
        traffic_data[988].size_bytes = 64;
        traffic_data[989].timestamp = 628;
        traffic_data[989].source_node = 9;
        traffic_data[989].dest_node = 3;
        traffic_data[989].packet_type = "CHI_READ";
        traffic_data[989].size_bytes = 64;
        traffic_data[990].timestamp = 628;
        traffic_data[990].source_node = 15;
        traffic_data[990].dest_node = 12;
        traffic_data[990].packet_type = "AXI_READ";
        traffic_data[990].size_bytes = 64;
        traffic_data[991].timestamp = 630;
        traffic_data[991].source_node = 6;
        traffic_data[991].dest_node = 9;
        traffic_data[991].packet_type = "CHI_READ";
        traffic_data[991].size_bytes = 64;
        traffic_data[992].timestamp = 630;
        traffic_data[992].source_node = 7;
        traffic_data[992].dest_node = 6;
        traffic_data[992].packet_type = "AXI_READ";
        traffic_data[992].size_bytes = 64;
        traffic_data[993].timestamp = 630;
        traffic_data[993].source_node = 14;
        traffic_data[993].dest_node = 1;
        traffic_data[993].packet_type = "AXI_READ";
        traffic_data[993].size_bytes = 64;
        traffic_data[994].timestamp = 631;
        traffic_data[994].source_node = 4;
        traffic_data[994].dest_node = 15;
        traffic_data[994].packet_type = "CHI_WRITE";
        traffic_data[994].size_bytes = 64;
        traffic_data[995].timestamp = 631;
        traffic_data[995].source_node = 15;
        traffic_data[995].dest_node = 10;
        traffic_data[995].packet_type = "CHI_READ";
        traffic_data[995].size_bytes = 64;
        traffic_data[996].timestamp = 632;
        traffic_data[996].source_node = 9;
        traffic_data[996].dest_node = 5;
        traffic_data[996].packet_type = "CHI_WRITE";
        traffic_data[996].size_bytes = 64;
        traffic_data[997].timestamp = 633;
        traffic_data[997].source_node = 12;
        traffic_data[997].dest_node = 2;
        traffic_data[997].packet_type = "CHI_READ";
        traffic_data[997].size_bytes = 64;
        traffic_data[998].timestamp = 635;
        traffic_data[998].source_node = 6;
        traffic_data[998].dest_node = 2;
        traffic_data[998].packet_type = "AXI_READ";
        traffic_data[998].size_bytes = 64;
        traffic_data[999].timestamp = 635;
        traffic_data[999].source_node = 15;
        traffic_data[999].dest_node = 8;
        traffic_data[999].packet_type = "CHI_READ";
        traffic_data[999].size_bytes = 64;
        traffic_data[1000].timestamp = 636;
        traffic_data[1000].source_node = 3;
        traffic_data[1000].dest_node = 7;
        traffic_data[1000].packet_type = "CHI_WRITE";
        traffic_data[1000].size_bytes = 64;
        traffic_data[1001].timestamp = 636;
        traffic_data[1001].source_node = 13;
        traffic_data[1001].dest_node = 10;
        traffic_data[1001].packet_type = "CHI_WRITE";
        traffic_data[1001].size_bytes = 64;
        traffic_data[1002].timestamp = 636;
        traffic_data[1002].source_node = 15;
        traffic_data[1002].dest_node = 4;
        traffic_data[1002].packet_type = "CHI_READ";
        traffic_data[1002].size_bytes = 64;
        traffic_data[1003].timestamp = 637;
        traffic_data[1003].source_node = 0;
        traffic_data[1003].dest_node = 14;
        traffic_data[1003].packet_type = "AXI_WRITE";
        traffic_data[1003].size_bytes = 64;
        traffic_data[1004].timestamp = 637;
        traffic_data[1004].source_node = 2;
        traffic_data[1004].dest_node = 9;
        traffic_data[1004].packet_type = "AXI_WRITE";
        traffic_data[1004].size_bytes = 64;
        traffic_data[1005].timestamp = 637;
        traffic_data[1005].source_node = 5;
        traffic_data[1005].dest_node = 10;
        traffic_data[1005].packet_type = "AXI_WRITE";
        traffic_data[1005].size_bytes = 64;
        traffic_data[1006].timestamp = 638;
        traffic_data[1006].source_node = 13;
        traffic_data[1006].dest_node = 14;
        traffic_data[1006].packet_type = "AXI_WRITE";
        traffic_data[1006].size_bytes = 64;
        traffic_data[1007].timestamp = 638;
        traffic_data[1007].source_node = 15;
        traffic_data[1007].dest_node = 6;
        traffic_data[1007].packet_type = "AXI_WRITE";
        traffic_data[1007].size_bytes = 64;
        traffic_data[1008].timestamp = 639;
        traffic_data[1008].source_node = 1;
        traffic_data[1008].dest_node = 15;
        traffic_data[1008].packet_type = "AXI_WRITE";
        traffic_data[1008].size_bytes = 64;
        traffic_data[1009].timestamp = 639;
        traffic_data[1009].source_node = 2;
        traffic_data[1009].dest_node = 1;
        traffic_data[1009].packet_type = "AXI_READ";
        traffic_data[1009].size_bytes = 64;
        traffic_data[1010].timestamp = 639;
        traffic_data[1010].source_node = 10;
        traffic_data[1010].dest_node = 7;
        traffic_data[1010].packet_type = "CHI_WRITE";
        traffic_data[1010].size_bytes = 64;
        traffic_data[1011].timestamp = 640;
        traffic_data[1011].source_node = 1;
        traffic_data[1011].dest_node = 8;
        traffic_data[1011].packet_type = "AXI_WRITE";
        traffic_data[1011].size_bytes = 64;
        traffic_data[1012].timestamp = 642;
        traffic_data[1012].source_node = 0;
        traffic_data[1012].dest_node = 11;
        traffic_data[1012].packet_type = "AXI_READ";
        traffic_data[1012].size_bytes = 64;
        traffic_data[1013].timestamp = 642;
        traffic_data[1013].source_node = 4;
        traffic_data[1013].dest_node = 8;
        traffic_data[1013].packet_type = "CHI_WRITE";
        traffic_data[1013].size_bytes = 64;
        traffic_data[1014].timestamp = 643;
        traffic_data[1014].source_node = 8;
        traffic_data[1014].dest_node = 14;
        traffic_data[1014].packet_type = "CHI_READ";
        traffic_data[1014].size_bytes = 64;
        traffic_data[1015].timestamp = 643;
        traffic_data[1015].source_node = 13;
        traffic_data[1015].dest_node = 8;
        traffic_data[1015].packet_type = "AXI_WRITE";
        traffic_data[1015].size_bytes = 64;
        traffic_data[1016].timestamp = 643;
        traffic_data[1016].source_node = 14;
        traffic_data[1016].dest_node = 7;
        traffic_data[1016].packet_type = "AXI_READ";
        traffic_data[1016].size_bytes = 64;
        traffic_data[1017].timestamp = 645;
        traffic_data[1017].source_node = 5;
        traffic_data[1017].dest_node = 9;
        traffic_data[1017].packet_type = "CHI_READ";
        traffic_data[1017].size_bytes = 64;
        traffic_data[1018].timestamp = 646;
        traffic_data[1018].source_node = 5;
        traffic_data[1018].dest_node = 7;
        traffic_data[1018].packet_type = "CHI_READ";
        traffic_data[1018].size_bytes = 64;
        traffic_data[1019].timestamp = 646;
        traffic_data[1019].source_node = 13;
        traffic_data[1019].dest_node = 11;
        traffic_data[1019].packet_type = "CHI_READ";
        traffic_data[1019].size_bytes = 64;
        traffic_data[1020].timestamp = 647;
        traffic_data[1020].source_node = 1;
        traffic_data[1020].dest_node = 13;
        traffic_data[1020].packet_type = "CHI_WRITE";
        traffic_data[1020].size_bytes = 64;
        traffic_data[1021].timestamp = 649;
        traffic_data[1021].source_node = 9;
        traffic_data[1021].dest_node = 14;
        traffic_data[1021].packet_type = "CHI_READ";
        traffic_data[1021].size_bytes = 64;
        traffic_data[1022].timestamp = 651;
        traffic_data[1022].source_node = 6;
        traffic_data[1022].dest_node = 1;
        traffic_data[1022].packet_type = "CHI_WRITE";
        traffic_data[1022].size_bytes = 64;
        traffic_data[1023].timestamp = 653;
        traffic_data[1023].source_node = 11;
        traffic_data[1023].dest_node = 9;
        traffic_data[1023].packet_type = "AXI_WRITE";
        traffic_data[1023].size_bytes = 64;
        traffic_data[1024].timestamp = 653;
        traffic_data[1024].source_node = 12;
        traffic_data[1024].dest_node = 5;
        traffic_data[1024].packet_type = "AXI_READ";
        traffic_data[1024].size_bytes = 64;
        traffic_data[1025].timestamp = 653;
        traffic_data[1025].source_node = 15;
        traffic_data[1025].dest_node = 7;
        traffic_data[1025].packet_type = "CHI_READ";
        traffic_data[1025].size_bytes = 64;
        traffic_data[1026].timestamp = 655;
        traffic_data[1026].source_node = 3;
        traffic_data[1026].dest_node = 6;
        traffic_data[1026].packet_type = "AXI_WRITE";
        traffic_data[1026].size_bytes = 64;
        traffic_data[1027].timestamp = 655;
        traffic_data[1027].source_node = 7;
        traffic_data[1027].dest_node = 6;
        traffic_data[1027].packet_type = "CHI_READ";
        traffic_data[1027].size_bytes = 64;
        traffic_data[1028].timestamp = 656;
        traffic_data[1028].source_node = 3;
        traffic_data[1028].dest_node = 4;
        traffic_data[1028].packet_type = "CHI_READ";
        traffic_data[1028].size_bytes = 64;
        traffic_data[1029].timestamp = 656;
        traffic_data[1029].source_node = 12;
        traffic_data[1029].dest_node = 9;
        traffic_data[1029].packet_type = "CHI_WRITE";
        traffic_data[1029].size_bytes = 64;
        traffic_data[1030].timestamp = 657;
        traffic_data[1030].source_node = 15;
        traffic_data[1030].dest_node = 3;
        traffic_data[1030].packet_type = "AXI_WRITE";
        traffic_data[1030].size_bytes = 64;
        traffic_data[1031].timestamp = 658;
        traffic_data[1031].source_node = 4;
        traffic_data[1031].dest_node = 3;
        traffic_data[1031].packet_type = "AXI_READ";
        traffic_data[1031].size_bytes = 64;
        traffic_data[1032].timestamp = 659;
        traffic_data[1032].source_node = 10;
        traffic_data[1032].dest_node = 12;
        traffic_data[1032].packet_type = "AXI_WRITE";
        traffic_data[1032].size_bytes = 64;
        traffic_data[1033].timestamp = 660;
        traffic_data[1033].source_node = 0;
        traffic_data[1033].dest_node = 15;
        traffic_data[1033].packet_type = "CHI_WRITE";
        traffic_data[1033].size_bytes = 64;
        traffic_data[1034].timestamp = 660;
        traffic_data[1034].source_node = 15;
        traffic_data[1034].dest_node = 2;
        traffic_data[1034].packet_type = "AXI_READ";
        traffic_data[1034].size_bytes = 64;
        traffic_data[1035].timestamp = 661;
        traffic_data[1035].source_node = 2;
        traffic_data[1035].dest_node = 6;
        traffic_data[1035].packet_type = "CHI_WRITE";
        traffic_data[1035].size_bytes = 64;
        traffic_data[1036].timestamp = 661;
        traffic_data[1036].source_node = 6;
        traffic_data[1036].dest_node = 12;
        traffic_data[1036].packet_type = "CHI_READ";
        traffic_data[1036].size_bytes = 64;
        traffic_data[1037].timestamp = 662;
        traffic_data[1037].source_node = 11;
        traffic_data[1037].dest_node = 9;
        traffic_data[1037].packet_type = "AXI_READ";
        traffic_data[1037].size_bytes = 64;
        traffic_data[1038].timestamp = 663;
        traffic_data[1038].source_node = 12;
        traffic_data[1038].dest_node = 6;
        traffic_data[1038].packet_type = "CHI_WRITE";
        traffic_data[1038].size_bytes = 64;
        traffic_data[1039].timestamp = 664;
        traffic_data[1039].source_node = 6;
        traffic_data[1039].dest_node = 4;
        traffic_data[1039].packet_type = "CHI_WRITE";
        traffic_data[1039].size_bytes = 64;
        traffic_data[1040].timestamp = 664;
        traffic_data[1040].source_node = 10;
        traffic_data[1040].dest_node = 7;
        traffic_data[1040].packet_type = "AXI_READ";
        traffic_data[1040].size_bytes = 64;
        traffic_data[1041].timestamp = 664;
        traffic_data[1041].source_node = 12;
        traffic_data[1041].dest_node = 9;
        traffic_data[1041].packet_type = "AXI_READ";
        traffic_data[1041].size_bytes = 64;
        traffic_data[1042].timestamp = 664;
        traffic_data[1042].source_node = 14;
        traffic_data[1042].dest_node = 5;
        traffic_data[1042].packet_type = "AXI_READ";
        traffic_data[1042].size_bytes = 64;
        traffic_data[1043].timestamp = 665;
        traffic_data[1043].source_node = 2;
        traffic_data[1043].dest_node = 7;
        traffic_data[1043].packet_type = "CHI_READ";
        traffic_data[1043].size_bytes = 64;
        traffic_data[1044].timestamp = 665;
        traffic_data[1044].source_node = 3;
        traffic_data[1044].dest_node = 15;
        traffic_data[1044].packet_type = "CHI_READ";
        traffic_data[1044].size_bytes = 64;
        traffic_data[1045].timestamp = 666;
        traffic_data[1045].source_node = 5;
        traffic_data[1045].dest_node = 0;
        traffic_data[1045].packet_type = "AXI_READ";
        traffic_data[1045].size_bytes = 64;
        traffic_data[1046].timestamp = 668;
        traffic_data[1046].source_node = 5;
        traffic_data[1046].dest_node = 9;
        traffic_data[1046].packet_type = "AXI_READ";
        traffic_data[1046].size_bytes = 64;
        traffic_data[1047].timestamp = 669;
        traffic_data[1047].source_node = 4;
        traffic_data[1047].dest_node = 0;
        traffic_data[1047].packet_type = "CHI_WRITE";
        traffic_data[1047].size_bytes = 64;
        traffic_data[1048].timestamp = 669;
        traffic_data[1048].source_node = 14;
        traffic_data[1048].dest_node = 1;
        traffic_data[1048].packet_type = "CHI_READ";
        traffic_data[1048].size_bytes = 64;
        traffic_data[1049].timestamp = 670;
        traffic_data[1049].source_node = 4;
        traffic_data[1049].dest_node = 0;
        traffic_data[1049].packet_type = "AXI_READ";
        traffic_data[1049].size_bytes = 64;
        traffic_data[1050].timestamp = 671;
        traffic_data[1050].source_node = 0;
        traffic_data[1050].dest_node = 4;
        traffic_data[1050].packet_type = "AXI_READ";
        traffic_data[1050].size_bytes = 64;
        traffic_data[1051].timestamp = 671;
        traffic_data[1051].source_node = 9;
        traffic_data[1051].dest_node = 6;
        traffic_data[1051].packet_type = "AXI_WRITE";
        traffic_data[1051].size_bytes = 64;
        traffic_data[1052].timestamp = 673;
        traffic_data[1052].source_node = 3;
        traffic_data[1052].dest_node = 14;
        traffic_data[1052].packet_type = "CHI_WRITE";
        traffic_data[1052].size_bytes = 64;
        traffic_data[1053].timestamp = 673;
        traffic_data[1053].source_node = 9;
        traffic_data[1053].dest_node = 12;
        traffic_data[1053].packet_type = "CHI_WRITE";
        traffic_data[1053].size_bytes = 64;
        traffic_data[1054].timestamp = 673;
        traffic_data[1054].source_node = 10;
        traffic_data[1054].dest_node = 13;
        traffic_data[1054].packet_type = "CHI_WRITE";
        traffic_data[1054].size_bytes = 64;
        traffic_data[1055].timestamp = 673;
        traffic_data[1055].source_node = 13;
        traffic_data[1055].dest_node = 1;
        traffic_data[1055].packet_type = "AXI_READ";
        traffic_data[1055].size_bytes = 64;
        traffic_data[1056].timestamp = 674;
        traffic_data[1056].source_node = 0;
        traffic_data[1056].dest_node = 9;
        traffic_data[1056].packet_type = "CHI_READ";
        traffic_data[1056].size_bytes = 64;
        traffic_data[1057].timestamp = 674;
        traffic_data[1057].source_node = 14;
        traffic_data[1057].dest_node = 13;
        traffic_data[1057].packet_type = "CHI_WRITE";
        traffic_data[1057].size_bytes = 64;
        traffic_data[1058].timestamp = 675;
        traffic_data[1058].source_node = 1;
        traffic_data[1058].dest_node = 8;
        traffic_data[1058].packet_type = "AXI_READ";
        traffic_data[1058].size_bytes = 64;
        traffic_data[1059].timestamp = 675;
        traffic_data[1059].source_node = 3;
        traffic_data[1059].dest_node = 7;
        traffic_data[1059].packet_type = "AXI_WRITE";
        traffic_data[1059].size_bytes = 64;
        traffic_data[1060].timestamp = 675;
        traffic_data[1060].source_node = 4;
        traffic_data[1060].dest_node = 12;
        traffic_data[1060].packet_type = "AXI_READ";
        traffic_data[1060].size_bytes = 64;
        traffic_data[1061].timestamp = 675;
        traffic_data[1061].source_node = 10;
        traffic_data[1061].dest_node = 15;
        traffic_data[1061].packet_type = "AXI_WRITE";
        traffic_data[1061].size_bytes = 64;
        traffic_data[1062].timestamp = 675;
        traffic_data[1062].source_node = 13;
        traffic_data[1062].dest_node = 0;
        traffic_data[1062].packet_type = "AXI_WRITE";
        traffic_data[1062].size_bytes = 64;
        traffic_data[1063].timestamp = 676;
        traffic_data[1063].source_node = 7;
        traffic_data[1063].dest_node = 2;
        traffic_data[1063].packet_type = "AXI_WRITE";
        traffic_data[1063].size_bytes = 64;
        traffic_data[1064].timestamp = 676;
        traffic_data[1064].source_node = 10;
        traffic_data[1064].dest_node = 7;
        traffic_data[1064].packet_type = "AXI_READ";
        traffic_data[1064].size_bytes = 64;
        traffic_data[1065].timestamp = 677;
        traffic_data[1065].source_node = 2;
        traffic_data[1065].dest_node = 9;
        traffic_data[1065].packet_type = "AXI_READ";
        traffic_data[1065].size_bytes = 64;
        traffic_data[1066].timestamp = 678;
        traffic_data[1066].source_node = 2;
        traffic_data[1066].dest_node = 11;
        traffic_data[1066].packet_type = "CHI_WRITE";
        traffic_data[1066].size_bytes = 64;
        traffic_data[1067].timestamp = 679;
        traffic_data[1067].source_node = 9;
        traffic_data[1067].dest_node = 13;
        traffic_data[1067].packet_type = "CHI_READ";
        traffic_data[1067].size_bytes = 64;
        traffic_data[1068].timestamp = 682;
        traffic_data[1068].source_node = 0;
        traffic_data[1068].dest_node = 4;
        traffic_data[1068].packet_type = "CHI_READ";
        traffic_data[1068].size_bytes = 64;
        traffic_data[1069].timestamp = 683;
        traffic_data[1069].source_node = 13;
        traffic_data[1069].dest_node = 0;
        traffic_data[1069].packet_type = "AXI_READ";
        traffic_data[1069].size_bytes = 64;
        traffic_data[1070].timestamp = 683;
        traffic_data[1070].source_node = 15;
        traffic_data[1070].dest_node = 14;
        traffic_data[1070].packet_type = "CHI_READ";
        traffic_data[1070].size_bytes = 64;
        traffic_data[1071].timestamp = 686;
        traffic_data[1071].source_node = 1;
        traffic_data[1071].dest_node = 12;
        traffic_data[1071].packet_type = "CHI_READ";
        traffic_data[1071].size_bytes = 64;
        traffic_data[1072].timestamp = 686;
        traffic_data[1072].source_node = 12;
        traffic_data[1072].dest_node = 2;
        traffic_data[1072].packet_type = "CHI_READ";
        traffic_data[1072].size_bytes = 64;
        traffic_data[1073].timestamp = 688;
        traffic_data[1073].source_node = 2;
        traffic_data[1073].dest_node = 6;
        traffic_data[1073].packet_type = "AXI_WRITE";
        traffic_data[1073].size_bytes = 64;
        traffic_data[1074].timestamp = 688;
        traffic_data[1074].source_node = 3;
        traffic_data[1074].dest_node = 4;
        traffic_data[1074].packet_type = "CHI_READ";
        traffic_data[1074].size_bytes = 64;
        traffic_data[1075].timestamp = 688;
        traffic_data[1075].source_node = 12;
        traffic_data[1075].dest_node = 14;
        traffic_data[1075].packet_type = "AXI_READ";
        traffic_data[1075].size_bytes = 64;
        traffic_data[1076].timestamp = 688;
        traffic_data[1076].source_node = 14;
        traffic_data[1076].dest_node = 6;
        traffic_data[1076].packet_type = "AXI_WRITE";
        traffic_data[1076].size_bytes = 64;
        traffic_data[1077].timestamp = 689;
        traffic_data[1077].source_node = 1;
        traffic_data[1077].dest_node = 11;
        traffic_data[1077].packet_type = "CHI_READ";
        traffic_data[1077].size_bytes = 64;
        traffic_data[1078].timestamp = 690;
        traffic_data[1078].source_node = 0;
        traffic_data[1078].dest_node = 11;
        traffic_data[1078].packet_type = "CHI_READ";
        traffic_data[1078].size_bytes = 64;
        traffic_data[1079].timestamp = 690;
        traffic_data[1079].source_node = 3;
        traffic_data[1079].dest_node = 2;
        traffic_data[1079].packet_type = "AXI_READ";
        traffic_data[1079].size_bytes = 64;
        traffic_data[1080].timestamp = 690;
        traffic_data[1080].source_node = 6;
        traffic_data[1080].dest_node = 10;
        traffic_data[1080].packet_type = "AXI_WRITE";
        traffic_data[1080].size_bytes = 64;
        traffic_data[1081].timestamp = 690;
        traffic_data[1081].source_node = 9;
        traffic_data[1081].dest_node = 0;
        traffic_data[1081].packet_type = "CHI_READ";
        traffic_data[1081].size_bytes = 64;
        traffic_data[1082].timestamp = 691;
        traffic_data[1082].source_node = 7;
        traffic_data[1082].dest_node = 1;
        traffic_data[1082].packet_type = "AXI_READ";
        traffic_data[1082].size_bytes = 64;
        traffic_data[1083].timestamp = 691;
        traffic_data[1083].source_node = 8;
        traffic_data[1083].dest_node = 13;
        traffic_data[1083].packet_type = "AXI_WRITE";
        traffic_data[1083].size_bytes = 64;
        traffic_data[1084].timestamp = 692;
        traffic_data[1084].source_node = 8;
        traffic_data[1084].dest_node = 3;
        traffic_data[1084].packet_type = "CHI_READ";
        traffic_data[1084].size_bytes = 64;
        traffic_data[1085].timestamp = 692;
        traffic_data[1085].source_node = 14;
        traffic_data[1085].dest_node = 2;
        traffic_data[1085].packet_type = "CHI_READ";
        traffic_data[1085].size_bytes = 64;
        traffic_data[1086].timestamp = 693;
        traffic_data[1086].source_node = 10;
        traffic_data[1086].dest_node = 15;
        traffic_data[1086].packet_type = "CHI_READ";
        traffic_data[1086].size_bytes = 64;
        traffic_data[1087].timestamp = 693;
        traffic_data[1087].source_node = 13;
        traffic_data[1087].dest_node = 7;
        traffic_data[1087].packet_type = "CHI_READ";
        traffic_data[1087].size_bytes = 64;
        traffic_data[1088].timestamp = 693;
        traffic_data[1088].source_node = 15;
        traffic_data[1088].dest_node = 12;
        traffic_data[1088].packet_type = "CHI_WRITE";
        traffic_data[1088].size_bytes = 64;
        traffic_data[1089].timestamp = 694;
        traffic_data[1089].source_node = 0;
        traffic_data[1089].dest_node = 13;
        traffic_data[1089].packet_type = "CHI_WRITE";
        traffic_data[1089].size_bytes = 64;
        traffic_data[1090].timestamp = 694;
        traffic_data[1090].source_node = 1;
        traffic_data[1090].dest_node = 12;
        traffic_data[1090].packet_type = "AXI_READ";
        traffic_data[1090].size_bytes = 64;
        traffic_data[1091].timestamp = 696;
        traffic_data[1091].source_node = 13;
        traffic_data[1091].dest_node = 7;
        traffic_data[1091].packet_type = "AXI_WRITE";
        traffic_data[1091].size_bytes = 64;
        traffic_data[1092].timestamp = 699;
        traffic_data[1092].source_node = 4;
        traffic_data[1092].dest_node = 6;
        traffic_data[1092].packet_type = "CHI_WRITE";
        traffic_data[1092].size_bytes = 64;
        traffic_data[1093].timestamp = 701;
        traffic_data[1093].source_node = 6;
        traffic_data[1093].dest_node = 7;
        traffic_data[1093].packet_type = "AXI_WRITE";
        traffic_data[1093].size_bytes = 64;
        traffic_data[1094].timestamp = 701;
        traffic_data[1094].source_node = 11;
        traffic_data[1094].dest_node = 3;
        traffic_data[1094].packet_type = "AXI_WRITE";
        traffic_data[1094].size_bytes = 64;
        traffic_data[1095].timestamp = 703;
        traffic_data[1095].source_node = 3;
        traffic_data[1095].dest_node = 5;
        traffic_data[1095].packet_type = "AXI_WRITE";
        traffic_data[1095].size_bytes = 64;
        traffic_data[1096].timestamp = 703;
        traffic_data[1096].source_node = 5;
        traffic_data[1096].dest_node = 11;
        traffic_data[1096].packet_type = "CHI_WRITE";
        traffic_data[1096].size_bytes = 64;
        traffic_data[1097].timestamp = 703;
        traffic_data[1097].source_node = 6;
        traffic_data[1097].dest_node = 8;
        traffic_data[1097].packet_type = "AXI_WRITE";
        traffic_data[1097].size_bytes = 64;
        traffic_data[1098].timestamp = 704;
        traffic_data[1098].source_node = 3;
        traffic_data[1098].dest_node = 0;
        traffic_data[1098].packet_type = "CHI_READ";
        traffic_data[1098].size_bytes = 64;
        traffic_data[1099].timestamp = 704;
        traffic_data[1099].source_node = 14;
        traffic_data[1099].dest_node = 4;
        traffic_data[1099].packet_type = "CHI_READ";
        traffic_data[1099].size_bytes = 64;
        traffic_data[1100].timestamp = 705;
        traffic_data[1100].source_node = 2;
        traffic_data[1100].dest_node = 12;
        traffic_data[1100].packet_type = "AXI_WRITE";
        traffic_data[1100].size_bytes = 64;
        traffic_data[1101].timestamp = 705;
        traffic_data[1101].source_node = 9;
        traffic_data[1101].dest_node = 5;
        traffic_data[1101].packet_type = "CHI_READ";
        traffic_data[1101].size_bytes = 64;
        traffic_data[1102].timestamp = 706;
        traffic_data[1102].source_node = 12;
        traffic_data[1102].dest_node = 14;
        traffic_data[1102].packet_type = "AXI_WRITE";
        traffic_data[1102].size_bytes = 64;
        traffic_data[1103].timestamp = 706;
        traffic_data[1103].source_node = 14;
        traffic_data[1103].dest_node = 12;
        traffic_data[1103].packet_type = "AXI_WRITE";
        traffic_data[1103].size_bytes = 64;
        traffic_data[1104].timestamp = 707;
        traffic_data[1104].source_node = 8;
        traffic_data[1104].dest_node = 12;
        traffic_data[1104].packet_type = "CHI_WRITE";
        traffic_data[1104].size_bytes = 64;
        traffic_data[1105].timestamp = 707;
        traffic_data[1105].source_node = 10;
        traffic_data[1105].dest_node = 9;
        traffic_data[1105].packet_type = "AXI_READ";
        traffic_data[1105].size_bytes = 64;
        traffic_data[1106].timestamp = 707;
        traffic_data[1106].source_node = 13;
        traffic_data[1106].dest_node = 11;
        traffic_data[1106].packet_type = "AXI_READ";
        traffic_data[1106].size_bytes = 64;
        traffic_data[1107].timestamp = 709;
        traffic_data[1107].source_node = 1;
        traffic_data[1107].dest_node = 10;
        traffic_data[1107].packet_type = "CHI_WRITE";
        traffic_data[1107].size_bytes = 64;
        traffic_data[1108].timestamp = 710;
        traffic_data[1108].source_node = 5;
        traffic_data[1108].dest_node = 0;
        traffic_data[1108].packet_type = "AXI_WRITE";
        traffic_data[1108].size_bytes = 64;
        traffic_data[1109].timestamp = 712;
        traffic_data[1109].source_node = 0;
        traffic_data[1109].dest_node = 4;
        traffic_data[1109].packet_type = "AXI_WRITE";
        traffic_data[1109].size_bytes = 64;
        traffic_data[1110].timestamp = 712;
        traffic_data[1110].source_node = 7;
        traffic_data[1110].dest_node = 1;
        traffic_data[1110].packet_type = "CHI_READ";
        traffic_data[1110].size_bytes = 64;
        traffic_data[1111].timestamp = 713;
        traffic_data[1111].source_node = 10;
        traffic_data[1111].dest_node = 9;
        traffic_data[1111].packet_type = "CHI_WRITE";
        traffic_data[1111].size_bytes = 64;
        traffic_data[1112].timestamp = 713;
        traffic_data[1112].source_node = 11;
        traffic_data[1112].dest_node = 12;
        traffic_data[1112].packet_type = "AXI_WRITE";
        traffic_data[1112].size_bytes = 64;
        traffic_data[1113].timestamp = 713;
        traffic_data[1113].source_node = 15;
        traffic_data[1113].dest_node = 6;
        traffic_data[1113].packet_type = "CHI_WRITE";
        traffic_data[1113].size_bytes = 64;
        traffic_data[1114].timestamp = 714;
        traffic_data[1114].source_node = 3;
        traffic_data[1114].dest_node = 1;
        traffic_data[1114].packet_type = "CHI_READ";
        traffic_data[1114].size_bytes = 64;
        traffic_data[1115].timestamp = 714;
        traffic_data[1115].source_node = 14;
        traffic_data[1115].dest_node = 9;
        traffic_data[1115].packet_type = "CHI_WRITE";
        traffic_data[1115].size_bytes = 64;
        traffic_data[1116].timestamp = 715;
        traffic_data[1116].source_node = 5;
        traffic_data[1116].dest_node = 6;
        traffic_data[1116].packet_type = "CHI_WRITE";
        traffic_data[1116].size_bytes = 64;
        traffic_data[1117].timestamp = 716;
        traffic_data[1117].source_node = 9;
        traffic_data[1117].dest_node = 4;
        traffic_data[1117].packet_type = "AXI_WRITE";
        traffic_data[1117].size_bytes = 64;
        traffic_data[1118].timestamp = 717;
        traffic_data[1118].source_node = 0;
        traffic_data[1118].dest_node = 9;
        traffic_data[1118].packet_type = "AXI_WRITE";
        traffic_data[1118].size_bytes = 64;
        traffic_data[1119].timestamp = 717;
        traffic_data[1119].source_node = 10;
        traffic_data[1119].dest_node = 6;
        traffic_data[1119].packet_type = "AXI_READ";
        traffic_data[1119].size_bytes = 64;
        traffic_data[1120].timestamp = 719;
        traffic_data[1120].source_node = 6;
        traffic_data[1120].dest_node = 13;
        traffic_data[1120].packet_type = "AXI_READ";
        traffic_data[1120].size_bytes = 64;
        traffic_data[1121].timestamp = 720;
        traffic_data[1121].source_node = 1;
        traffic_data[1121].dest_node = 5;
        traffic_data[1121].packet_type = "AXI_READ";
        traffic_data[1121].size_bytes = 64;
        traffic_data[1122].timestamp = 720;
        traffic_data[1122].source_node = 5;
        traffic_data[1122].dest_node = 8;
        traffic_data[1122].packet_type = "AXI_READ";
        traffic_data[1122].size_bytes = 64;
        traffic_data[1123].timestamp = 721;
        traffic_data[1123].source_node = 1;
        traffic_data[1123].dest_node = 8;
        traffic_data[1123].packet_type = "AXI_READ";
        traffic_data[1123].size_bytes = 64;
        traffic_data[1124].timestamp = 722;
        traffic_data[1124].source_node = 2;
        traffic_data[1124].dest_node = 5;
        traffic_data[1124].packet_type = "AXI_READ";
        traffic_data[1124].size_bytes = 64;
        traffic_data[1125].timestamp = 722;
        traffic_data[1125].source_node = 3;
        traffic_data[1125].dest_node = 12;
        traffic_data[1125].packet_type = "AXI_READ";
        traffic_data[1125].size_bytes = 64;
        traffic_data[1126].timestamp = 722;
        traffic_data[1126].source_node = 8;
        traffic_data[1126].dest_node = 4;
        traffic_data[1126].packet_type = "CHI_WRITE";
        traffic_data[1126].size_bytes = 64;
        traffic_data[1127].timestamp = 722;
        traffic_data[1127].source_node = 11;
        traffic_data[1127].dest_node = 2;
        traffic_data[1127].packet_type = "AXI_READ";
        traffic_data[1127].size_bytes = 64;
        traffic_data[1128].timestamp = 723;
        traffic_data[1128].source_node = 4;
        traffic_data[1128].dest_node = 10;
        traffic_data[1128].packet_type = "AXI_READ";
        traffic_data[1128].size_bytes = 64;
        traffic_data[1129].timestamp = 724;
        traffic_data[1129].source_node = 1;
        traffic_data[1129].dest_node = 13;
        traffic_data[1129].packet_type = "AXI_WRITE";
        traffic_data[1129].size_bytes = 64;
        traffic_data[1130].timestamp = 724;
        traffic_data[1130].source_node = 3;
        traffic_data[1130].dest_node = 2;
        traffic_data[1130].packet_type = "AXI_WRITE";
        traffic_data[1130].size_bytes = 64;
        traffic_data[1131].timestamp = 725;
        traffic_data[1131].source_node = 3;
        traffic_data[1131].dest_node = 9;
        traffic_data[1131].packet_type = "CHI_READ";
        traffic_data[1131].size_bytes = 64;
        traffic_data[1132].timestamp = 725;
        traffic_data[1132].source_node = 10;
        traffic_data[1132].dest_node = 4;
        traffic_data[1132].packet_type = "CHI_READ";
        traffic_data[1132].size_bytes = 64;
        traffic_data[1133].timestamp = 726;
        traffic_data[1133].source_node = 0;
        traffic_data[1133].dest_node = 2;
        traffic_data[1133].packet_type = "AXI_WRITE";
        traffic_data[1133].size_bytes = 64;
        traffic_data[1134].timestamp = 726;
        traffic_data[1134].source_node = 6;
        traffic_data[1134].dest_node = 13;
        traffic_data[1134].packet_type = "AXI_WRITE";
        traffic_data[1134].size_bytes = 64;
        traffic_data[1135].timestamp = 726;
        traffic_data[1135].source_node = 9;
        traffic_data[1135].dest_node = 3;
        traffic_data[1135].packet_type = "AXI_WRITE";
        traffic_data[1135].size_bytes = 64;
        traffic_data[1136].timestamp = 726;
        traffic_data[1136].source_node = 15;
        traffic_data[1136].dest_node = 8;
        traffic_data[1136].packet_type = "CHI_READ";
        traffic_data[1136].size_bytes = 64;
        traffic_data[1137].timestamp = 727;
        traffic_data[1137].source_node = 1;
        traffic_data[1137].dest_node = 15;
        traffic_data[1137].packet_type = "AXI_WRITE";
        traffic_data[1137].size_bytes = 64;
        traffic_data[1138].timestamp = 727;
        traffic_data[1138].source_node = 13;
        traffic_data[1138].dest_node = 10;
        traffic_data[1138].packet_type = "AXI_WRITE";
        traffic_data[1138].size_bytes = 64;
        traffic_data[1139].timestamp = 728;
        traffic_data[1139].source_node = 3;
        traffic_data[1139].dest_node = 2;
        traffic_data[1139].packet_type = "AXI_WRITE";
        traffic_data[1139].size_bytes = 64;
        traffic_data[1140].timestamp = 728;
        traffic_data[1140].source_node = 11;
        traffic_data[1140].dest_node = 5;
        traffic_data[1140].packet_type = "CHI_WRITE";
        traffic_data[1140].size_bytes = 64;
        traffic_data[1141].timestamp = 728;
        traffic_data[1141].source_node = 12;
        traffic_data[1141].dest_node = 10;
        traffic_data[1141].packet_type = "CHI_READ";
        traffic_data[1141].size_bytes = 64;
        traffic_data[1142].timestamp = 729;
        traffic_data[1142].source_node = 12;
        traffic_data[1142].dest_node = 1;
        traffic_data[1142].packet_type = "AXI_READ";
        traffic_data[1142].size_bytes = 64;
        traffic_data[1143].timestamp = 730;
        traffic_data[1143].source_node = 0;
        traffic_data[1143].dest_node = 5;
        traffic_data[1143].packet_type = "CHI_WRITE";
        traffic_data[1143].size_bytes = 64;
        traffic_data[1144].timestamp = 731;
        traffic_data[1144].source_node = 8;
        traffic_data[1144].dest_node = 11;
        traffic_data[1144].packet_type = "CHI_READ";
        traffic_data[1144].size_bytes = 64;
        traffic_data[1145].timestamp = 734;
        traffic_data[1145].source_node = 4;
        traffic_data[1145].dest_node = 1;
        traffic_data[1145].packet_type = "CHI_WRITE";
        traffic_data[1145].size_bytes = 64;
        traffic_data[1146].timestamp = 734;
        traffic_data[1146].source_node = 7;
        traffic_data[1146].dest_node = 3;
        traffic_data[1146].packet_type = "CHI_READ";
        traffic_data[1146].size_bytes = 64;
        traffic_data[1147].timestamp = 734;
        traffic_data[1147].source_node = 15;
        traffic_data[1147].dest_node = 6;
        traffic_data[1147].packet_type = "CHI_WRITE";
        traffic_data[1147].size_bytes = 64;
        traffic_data[1148].timestamp = 735;
        traffic_data[1148].source_node = 7;
        traffic_data[1148].dest_node = 14;
        traffic_data[1148].packet_type = "AXI_READ";
        traffic_data[1148].size_bytes = 64;
        traffic_data[1149].timestamp = 736;
        traffic_data[1149].source_node = 1;
        traffic_data[1149].dest_node = 6;
        traffic_data[1149].packet_type = "CHI_READ";
        traffic_data[1149].size_bytes = 64;
        traffic_data[1150].timestamp = 736;
        traffic_data[1150].source_node = 10;
        traffic_data[1150].dest_node = 9;
        traffic_data[1150].packet_type = "CHI_READ";
        traffic_data[1150].size_bytes = 64;
        traffic_data[1151].timestamp = 737;
        traffic_data[1151].source_node = 0;
        traffic_data[1151].dest_node = 3;
        traffic_data[1151].packet_type = "AXI_READ";
        traffic_data[1151].size_bytes = 64;
        traffic_data[1152].timestamp = 737;
        traffic_data[1152].source_node = 13;
        traffic_data[1152].dest_node = 10;
        traffic_data[1152].packet_type = "CHI_READ";
        traffic_data[1152].size_bytes = 64;
        traffic_data[1153].timestamp = 738;
        traffic_data[1153].source_node = 10;
        traffic_data[1153].dest_node = 13;
        traffic_data[1153].packet_type = "CHI_READ";
        traffic_data[1153].size_bytes = 64;
        traffic_data[1154].timestamp = 739;
        traffic_data[1154].source_node = 0;
        traffic_data[1154].dest_node = 9;
        traffic_data[1154].packet_type = "CHI_WRITE";
        traffic_data[1154].size_bytes = 64;
        traffic_data[1155].timestamp = 740;
        traffic_data[1155].source_node = 1;
        traffic_data[1155].dest_node = 15;
        traffic_data[1155].packet_type = "AXI_WRITE";
        traffic_data[1155].size_bytes = 64;
        traffic_data[1156].timestamp = 740;
        traffic_data[1156].source_node = 3;
        traffic_data[1156].dest_node = 12;
        traffic_data[1156].packet_type = "AXI_READ";
        traffic_data[1156].size_bytes = 64;
        traffic_data[1157].timestamp = 740;
        traffic_data[1157].source_node = 10;
        traffic_data[1157].dest_node = 4;
        traffic_data[1157].packet_type = "CHI_READ";
        traffic_data[1157].size_bytes = 64;
        traffic_data[1158].timestamp = 741;
        traffic_data[1158].source_node = 8;
        traffic_data[1158].dest_node = 15;
        traffic_data[1158].packet_type = "AXI_WRITE";
        traffic_data[1158].size_bytes = 64;
        traffic_data[1159].timestamp = 741;
        traffic_data[1159].source_node = 9;
        traffic_data[1159].dest_node = 12;
        traffic_data[1159].packet_type = "AXI_READ";
        traffic_data[1159].size_bytes = 64;
        traffic_data[1160].timestamp = 742;
        traffic_data[1160].source_node = 4;
        traffic_data[1160].dest_node = 14;
        traffic_data[1160].packet_type = "AXI_READ";
        traffic_data[1160].size_bytes = 64;
        traffic_data[1161].timestamp = 742;
        traffic_data[1161].source_node = 15;
        traffic_data[1161].dest_node = 3;
        traffic_data[1161].packet_type = "AXI_READ";
        traffic_data[1161].size_bytes = 64;
        traffic_data[1162].timestamp = 743;
        traffic_data[1162].source_node = 0;
        traffic_data[1162].dest_node = 2;
        traffic_data[1162].packet_type = "CHI_READ";
        traffic_data[1162].size_bytes = 64;
        traffic_data[1163].timestamp = 743;
        traffic_data[1163].source_node = 10;
        traffic_data[1163].dest_node = 14;
        traffic_data[1163].packet_type = "AXI_WRITE";
        traffic_data[1163].size_bytes = 64;
        traffic_data[1164].timestamp = 743;
        traffic_data[1164].source_node = 13;
        traffic_data[1164].dest_node = 8;
        traffic_data[1164].packet_type = "AXI_READ";
        traffic_data[1164].size_bytes = 64;
        traffic_data[1165].timestamp = 744;
        traffic_data[1165].source_node = 12;
        traffic_data[1165].dest_node = 6;
        traffic_data[1165].packet_type = "AXI_WRITE";
        traffic_data[1165].size_bytes = 64;
        traffic_data[1166].timestamp = 744;
        traffic_data[1166].source_node = 13;
        traffic_data[1166].dest_node = 7;
        traffic_data[1166].packet_type = "CHI_WRITE";
        traffic_data[1166].size_bytes = 64;
        traffic_data[1167].timestamp = 746;
        traffic_data[1167].source_node = 9;
        traffic_data[1167].dest_node = 6;
        traffic_data[1167].packet_type = "AXI_WRITE";
        traffic_data[1167].size_bytes = 64;
        traffic_data[1168].timestamp = 748;
        traffic_data[1168].source_node = 3;
        traffic_data[1168].dest_node = 5;
        traffic_data[1168].packet_type = "CHI_READ";
        traffic_data[1168].size_bytes = 64;
        traffic_data[1169].timestamp = 748;
        traffic_data[1169].source_node = 6;
        traffic_data[1169].dest_node = 14;
        traffic_data[1169].packet_type = "CHI_WRITE";
        traffic_data[1169].size_bytes = 64;
        traffic_data[1170].timestamp = 748;
        traffic_data[1170].source_node = 7;
        traffic_data[1170].dest_node = 5;
        traffic_data[1170].packet_type = "AXI_WRITE";
        traffic_data[1170].size_bytes = 64;
        traffic_data[1171].timestamp = 748;
        traffic_data[1171].source_node = 10;
        traffic_data[1171].dest_node = 1;
        traffic_data[1171].packet_type = "AXI_WRITE";
        traffic_data[1171].size_bytes = 64;
        traffic_data[1172].timestamp = 748;
        traffic_data[1172].source_node = 13;
        traffic_data[1172].dest_node = 8;
        traffic_data[1172].packet_type = "AXI_WRITE";
        traffic_data[1172].size_bytes = 64;
        traffic_data[1173].timestamp = 750;
        traffic_data[1173].source_node = 13;
        traffic_data[1173].dest_node = 0;
        traffic_data[1173].packet_type = "AXI_WRITE";
        traffic_data[1173].size_bytes = 64;
        traffic_data[1174].timestamp = 751;
        traffic_data[1174].source_node = 6;
        traffic_data[1174].dest_node = 1;
        traffic_data[1174].packet_type = "AXI_WRITE";
        traffic_data[1174].size_bytes = 64;
        traffic_data[1175].timestamp = 751;
        traffic_data[1175].source_node = 10;
        traffic_data[1175].dest_node = 7;
        traffic_data[1175].packet_type = "AXI_WRITE";
        traffic_data[1175].size_bytes = 64;
        traffic_data[1176].timestamp = 751;
        traffic_data[1176].source_node = 13;
        traffic_data[1176].dest_node = 7;
        traffic_data[1176].packet_type = "CHI_READ";
        traffic_data[1176].size_bytes = 64;
        traffic_data[1177].timestamp = 753;
        traffic_data[1177].source_node = 7;
        traffic_data[1177].dest_node = 10;
        traffic_data[1177].packet_type = "CHI_READ";
        traffic_data[1177].size_bytes = 64;
        traffic_data[1178].timestamp = 754;
        traffic_data[1178].source_node = 1;
        traffic_data[1178].dest_node = 9;
        traffic_data[1178].packet_type = "CHI_READ";
        traffic_data[1178].size_bytes = 64;
        traffic_data[1179].timestamp = 754;
        traffic_data[1179].source_node = 12;
        traffic_data[1179].dest_node = 6;
        traffic_data[1179].packet_type = "CHI_WRITE";
        traffic_data[1179].size_bytes = 64;
        traffic_data[1180].timestamp = 754;
        traffic_data[1180].source_node = 15;
        traffic_data[1180].dest_node = 5;
        traffic_data[1180].packet_type = "AXI_READ";
        traffic_data[1180].size_bytes = 64;
        traffic_data[1181].timestamp = 755;
        traffic_data[1181].source_node = 15;
        traffic_data[1181].dest_node = 11;
        traffic_data[1181].packet_type = "AXI_READ";
        traffic_data[1181].size_bytes = 64;
        traffic_data[1182].timestamp = 756;
        traffic_data[1182].source_node = 7;
        traffic_data[1182].dest_node = 8;
        traffic_data[1182].packet_type = "AXI_WRITE";
        traffic_data[1182].size_bytes = 64;
        traffic_data[1183].timestamp = 756;
        traffic_data[1183].source_node = 8;
        traffic_data[1183].dest_node = 4;
        traffic_data[1183].packet_type = "CHI_READ";
        traffic_data[1183].size_bytes = 64;
        traffic_data[1184].timestamp = 756;
        traffic_data[1184].source_node = 13;
        traffic_data[1184].dest_node = 2;
        traffic_data[1184].packet_type = "CHI_READ";
        traffic_data[1184].size_bytes = 64;
        traffic_data[1185].timestamp = 756;
        traffic_data[1185].source_node = 15;
        traffic_data[1185].dest_node = 9;
        traffic_data[1185].packet_type = "AXI_READ";
        traffic_data[1185].size_bytes = 64;
        traffic_data[1186].timestamp = 757;
        traffic_data[1186].source_node = 13;
        traffic_data[1186].dest_node = 9;
        traffic_data[1186].packet_type = "CHI_READ";
        traffic_data[1186].size_bytes = 64;
        traffic_data[1187].timestamp = 759;
        traffic_data[1187].source_node = 5;
        traffic_data[1187].dest_node = 0;
        traffic_data[1187].packet_type = "AXI_READ";
        traffic_data[1187].size_bytes = 64;
        traffic_data[1188].timestamp = 760;
        traffic_data[1188].source_node = 11;
        traffic_data[1188].dest_node = 14;
        traffic_data[1188].packet_type = "CHI_READ";
        traffic_data[1188].size_bytes = 64;
        traffic_data[1189].timestamp = 761;
        traffic_data[1189].source_node = 14;
        traffic_data[1189].dest_node = 15;
        traffic_data[1189].packet_type = "CHI_READ";
        traffic_data[1189].size_bytes = 64;
        traffic_data[1190].timestamp = 762;
        traffic_data[1190].source_node = 12;
        traffic_data[1190].dest_node = 7;
        traffic_data[1190].packet_type = "AXI_WRITE";
        traffic_data[1190].size_bytes = 64;
        traffic_data[1191].timestamp = 763;
        traffic_data[1191].source_node = 15;
        traffic_data[1191].dest_node = 5;
        traffic_data[1191].packet_type = "AXI_READ";
        traffic_data[1191].size_bytes = 64;
        traffic_data[1192].timestamp = 764;
        traffic_data[1192].source_node = 14;
        traffic_data[1192].dest_node = 3;
        traffic_data[1192].packet_type = "CHI_READ";
        traffic_data[1192].size_bytes = 64;
        traffic_data[1193].timestamp = 765;
        traffic_data[1193].source_node = 0;
        traffic_data[1193].dest_node = 4;
        traffic_data[1193].packet_type = "AXI_READ";
        traffic_data[1193].size_bytes = 64;
        traffic_data[1194].timestamp = 765;
        traffic_data[1194].source_node = 4;
        traffic_data[1194].dest_node = 0;
        traffic_data[1194].packet_type = "AXI_READ";
        traffic_data[1194].size_bytes = 64;
        traffic_data[1195].timestamp = 766;
        traffic_data[1195].source_node = 0;
        traffic_data[1195].dest_node = 10;
        traffic_data[1195].packet_type = "AXI_WRITE";
        traffic_data[1195].size_bytes = 64;
        traffic_data[1196].timestamp = 766;
        traffic_data[1196].source_node = 10;
        traffic_data[1196].dest_node = 6;
        traffic_data[1196].packet_type = "AXI_READ";
        traffic_data[1196].size_bytes = 64;
        traffic_data[1197].timestamp = 766;
        traffic_data[1197].source_node = 14;
        traffic_data[1197].dest_node = 15;
        traffic_data[1197].packet_type = "CHI_READ";
        traffic_data[1197].size_bytes = 64;
        traffic_data[1198].timestamp = 767;
        traffic_data[1198].source_node = 11;
        traffic_data[1198].dest_node = 2;
        traffic_data[1198].packet_type = "AXI_READ";
        traffic_data[1198].size_bytes = 64;
        traffic_data[1199].timestamp = 767;
        traffic_data[1199].source_node = 13;
        traffic_data[1199].dest_node = 3;
        traffic_data[1199].packet_type = "AXI_READ";
        traffic_data[1199].size_bytes = 64;
        traffic_data[1200].timestamp = 768;
        traffic_data[1200].source_node = 11;
        traffic_data[1200].dest_node = 13;
        traffic_data[1200].packet_type = "AXI_READ";
        traffic_data[1200].size_bytes = 64;
        traffic_data[1201].timestamp = 770;
        traffic_data[1201].source_node = 9;
        traffic_data[1201].dest_node = 12;
        traffic_data[1201].packet_type = "AXI_WRITE";
        traffic_data[1201].size_bytes = 64;
        traffic_data[1202].timestamp = 771;
        traffic_data[1202].source_node = 2;
        traffic_data[1202].dest_node = 4;
        traffic_data[1202].packet_type = "AXI_READ";
        traffic_data[1202].size_bytes = 64;
        traffic_data[1203].timestamp = 771;
        traffic_data[1203].source_node = 4;
        traffic_data[1203].dest_node = 11;
        traffic_data[1203].packet_type = "CHI_READ";
        traffic_data[1203].size_bytes = 64;
        traffic_data[1204].timestamp = 771;
        traffic_data[1204].source_node = 10;
        traffic_data[1204].dest_node = 14;
        traffic_data[1204].packet_type = "AXI_READ";
        traffic_data[1204].size_bytes = 64;
        traffic_data[1205].timestamp = 772;
        traffic_data[1205].source_node = 4;
        traffic_data[1205].dest_node = 14;
        traffic_data[1205].packet_type = "CHI_READ";
        traffic_data[1205].size_bytes = 64;
        traffic_data[1206].timestamp = 772;
        traffic_data[1206].source_node = 8;
        traffic_data[1206].dest_node = 1;
        traffic_data[1206].packet_type = "AXI_READ";
        traffic_data[1206].size_bytes = 64;
        traffic_data[1207].timestamp = 773;
        traffic_data[1207].source_node = 7;
        traffic_data[1207].dest_node = 4;
        traffic_data[1207].packet_type = "CHI_READ";
        traffic_data[1207].size_bytes = 64;
        traffic_data[1208].timestamp = 773;
        traffic_data[1208].source_node = 9;
        traffic_data[1208].dest_node = 2;
        traffic_data[1208].packet_type = "AXI_READ";
        traffic_data[1208].size_bytes = 64;
        traffic_data[1209].timestamp = 773;
        traffic_data[1209].source_node = 11;
        traffic_data[1209].dest_node = 4;
        traffic_data[1209].packet_type = "CHI_READ";
        traffic_data[1209].size_bytes = 64;
        traffic_data[1210].timestamp = 774;
        traffic_data[1210].source_node = 0;
        traffic_data[1210].dest_node = 1;
        traffic_data[1210].packet_type = "CHI_READ";
        traffic_data[1210].size_bytes = 64;
        traffic_data[1211].timestamp = 774;
        traffic_data[1211].source_node = 5;
        traffic_data[1211].dest_node = 12;
        traffic_data[1211].packet_type = "CHI_READ";
        traffic_data[1211].size_bytes = 64;
        traffic_data[1212].timestamp = 774;
        traffic_data[1212].source_node = 13;
        traffic_data[1212].dest_node = 5;
        traffic_data[1212].packet_type = "CHI_READ";
        traffic_data[1212].size_bytes = 64;
        traffic_data[1213].timestamp = 775;
        traffic_data[1213].source_node = 0;
        traffic_data[1213].dest_node = 10;
        traffic_data[1213].packet_type = "AXI_READ";
        traffic_data[1213].size_bytes = 64;
        traffic_data[1214].timestamp = 775;
        traffic_data[1214].source_node = 10;
        traffic_data[1214].dest_node = 2;
        traffic_data[1214].packet_type = "AXI_WRITE";
        traffic_data[1214].size_bytes = 64;
        traffic_data[1215].timestamp = 775;
        traffic_data[1215].source_node = 15;
        traffic_data[1215].dest_node = 3;
        traffic_data[1215].packet_type = "AXI_WRITE";
        traffic_data[1215].size_bytes = 64;
        traffic_data[1216].timestamp = 776;
        traffic_data[1216].source_node = 5;
        traffic_data[1216].dest_node = 9;
        traffic_data[1216].packet_type = "CHI_READ";
        traffic_data[1216].size_bytes = 64;
        traffic_data[1217].timestamp = 777;
        traffic_data[1217].source_node = 10;
        traffic_data[1217].dest_node = 1;
        traffic_data[1217].packet_type = "CHI_WRITE";
        traffic_data[1217].size_bytes = 64;
        traffic_data[1218].timestamp = 778;
        traffic_data[1218].source_node = 6;
        traffic_data[1218].dest_node = 1;
        traffic_data[1218].packet_type = "CHI_WRITE";
        traffic_data[1218].size_bytes = 64;
        traffic_data[1219].timestamp = 778;
        traffic_data[1219].source_node = 14;
        traffic_data[1219].dest_node = 1;
        traffic_data[1219].packet_type = "CHI_READ";
        traffic_data[1219].size_bytes = 64;
        traffic_data[1220].timestamp = 781;
        traffic_data[1220].source_node = 2;
        traffic_data[1220].dest_node = 8;
        traffic_data[1220].packet_type = "CHI_READ";
        traffic_data[1220].size_bytes = 64;
        traffic_data[1221].timestamp = 782;
        traffic_data[1221].source_node = 7;
        traffic_data[1221].dest_node = 14;
        traffic_data[1221].packet_type = "CHI_READ";
        traffic_data[1221].size_bytes = 64;
        traffic_data[1222].timestamp = 782;
        traffic_data[1222].source_node = 9;
        traffic_data[1222].dest_node = 10;
        traffic_data[1222].packet_type = "AXI_READ";
        traffic_data[1222].size_bytes = 64;
        traffic_data[1223].timestamp = 783;
        traffic_data[1223].source_node = 7;
        traffic_data[1223].dest_node = 13;
        traffic_data[1223].packet_type = "CHI_WRITE";
        traffic_data[1223].size_bytes = 64;
        traffic_data[1224].timestamp = 783;
        traffic_data[1224].source_node = 9;
        traffic_data[1224].dest_node = 3;
        traffic_data[1224].packet_type = "AXI_WRITE";
        traffic_data[1224].size_bytes = 64;
        traffic_data[1225].timestamp = 785;
        traffic_data[1225].source_node = 8;
        traffic_data[1225].dest_node = 11;
        traffic_data[1225].packet_type = "CHI_WRITE";
        traffic_data[1225].size_bytes = 64;
        traffic_data[1226].timestamp = 785;
        traffic_data[1226].source_node = 13;
        traffic_data[1226].dest_node = 0;
        traffic_data[1226].packet_type = "CHI_WRITE";
        traffic_data[1226].size_bytes = 64;
        traffic_data[1227].timestamp = 786;
        traffic_data[1227].source_node = 11;
        traffic_data[1227].dest_node = 12;
        traffic_data[1227].packet_type = "CHI_READ";
        traffic_data[1227].size_bytes = 64;
        traffic_data[1228].timestamp = 786;
        traffic_data[1228].source_node = 15;
        traffic_data[1228].dest_node = 13;
        traffic_data[1228].packet_type = "CHI_WRITE";
        traffic_data[1228].size_bytes = 64;
        traffic_data[1229].timestamp = 787;
        traffic_data[1229].source_node = 4;
        traffic_data[1229].dest_node = 10;
        traffic_data[1229].packet_type = "AXI_WRITE";
        traffic_data[1229].size_bytes = 64;
        traffic_data[1230].timestamp = 787;
        traffic_data[1230].source_node = 12;
        traffic_data[1230].dest_node = 1;
        traffic_data[1230].packet_type = "AXI_READ";
        traffic_data[1230].size_bytes = 64;
        traffic_data[1231].timestamp = 788;
        traffic_data[1231].source_node = 1;
        traffic_data[1231].dest_node = 3;
        traffic_data[1231].packet_type = "AXI_WRITE";
        traffic_data[1231].size_bytes = 64;
        traffic_data[1232].timestamp = 788;
        traffic_data[1232].source_node = 5;
        traffic_data[1232].dest_node = 8;
        traffic_data[1232].packet_type = "AXI_WRITE";
        traffic_data[1232].size_bytes = 64;
        traffic_data[1233].timestamp = 788;
        traffic_data[1233].source_node = 7;
        traffic_data[1233].dest_node = 12;
        traffic_data[1233].packet_type = "AXI_WRITE";
        traffic_data[1233].size_bytes = 64;
        traffic_data[1234].timestamp = 789;
        traffic_data[1234].source_node = 2;
        traffic_data[1234].dest_node = 3;
        traffic_data[1234].packet_type = "CHI_WRITE";
        traffic_data[1234].size_bytes = 64;
        traffic_data[1235].timestamp = 791;
        traffic_data[1235].source_node = 1;
        traffic_data[1235].dest_node = 7;
        traffic_data[1235].packet_type = "CHI_READ";
        traffic_data[1235].size_bytes = 64;
        traffic_data[1236].timestamp = 793;
        traffic_data[1236].source_node = 10;
        traffic_data[1236].dest_node = 12;
        traffic_data[1236].packet_type = "AXI_READ";
        traffic_data[1236].size_bytes = 64;
        traffic_data[1237].timestamp = 794;
        traffic_data[1237].source_node = 0;
        traffic_data[1237].dest_node = 13;
        traffic_data[1237].packet_type = "AXI_READ";
        traffic_data[1237].size_bytes = 64;
        traffic_data[1238].timestamp = 794;
        traffic_data[1238].source_node = 6;
        traffic_data[1238].dest_node = 2;
        traffic_data[1238].packet_type = "AXI_READ";
        traffic_data[1238].size_bytes = 64;
        traffic_data[1239].timestamp = 794;
        traffic_data[1239].source_node = 7;
        traffic_data[1239].dest_node = 3;
        traffic_data[1239].packet_type = "CHI_WRITE";
        traffic_data[1239].size_bytes = 64;
        traffic_data[1240].timestamp = 794;
        traffic_data[1240].source_node = 9;
        traffic_data[1240].dest_node = 13;
        traffic_data[1240].packet_type = "CHI_READ";
        traffic_data[1240].size_bytes = 64;
        traffic_data[1241].timestamp = 794;
        traffic_data[1241].source_node = 10;
        traffic_data[1241].dest_node = 11;
        traffic_data[1241].packet_type = "AXI_READ";
        traffic_data[1241].size_bytes = 64;
        traffic_data[1242].timestamp = 795;
        traffic_data[1242].source_node = 15;
        traffic_data[1242].dest_node = 6;
        traffic_data[1242].packet_type = "CHI_WRITE";
        traffic_data[1242].size_bytes = 64;
        traffic_data[1243].timestamp = 796;
        traffic_data[1243].source_node = 0;
        traffic_data[1243].dest_node = 7;
        traffic_data[1243].packet_type = "CHI_WRITE";
        traffic_data[1243].size_bytes = 64;
        traffic_data[1244].timestamp = 796;
        traffic_data[1244].source_node = 1;
        traffic_data[1244].dest_node = 10;
        traffic_data[1244].packet_type = "AXI_READ";
        traffic_data[1244].size_bytes = 64;
        traffic_data[1245].timestamp = 796;
        traffic_data[1245].source_node = 2;
        traffic_data[1245].dest_node = 5;
        traffic_data[1245].packet_type = "AXI_WRITE";
        traffic_data[1245].size_bytes = 64;
        traffic_data[1246].timestamp = 796;
        traffic_data[1246].source_node = 5;
        traffic_data[1246].dest_node = 12;
        traffic_data[1246].packet_type = "CHI_READ";
        traffic_data[1246].size_bytes = 64;
        traffic_data[1247].timestamp = 797;
        traffic_data[1247].source_node = 3;
        traffic_data[1247].dest_node = 12;
        traffic_data[1247].packet_type = "AXI_READ";
        traffic_data[1247].size_bytes = 64;
        traffic_data[1248].timestamp = 797;
        traffic_data[1248].source_node = 5;
        traffic_data[1248].dest_node = 3;
        traffic_data[1248].packet_type = "AXI_WRITE";
        traffic_data[1248].size_bytes = 64;
        traffic_data[1249].timestamp = 797;
        traffic_data[1249].source_node = 11;
        traffic_data[1249].dest_node = 9;
        traffic_data[1249].packet_type = "AXI_WRITE";
        traffic_data[1249].size_bytes = 64;
        traffic_data[1250].timestamp = 797;
        traffic_data[1250].source_node = 13;
        traffic_data[1250].dest_node = 12;
        traffic_data[1250].packet_type = "AXI_READ";
        traffic_data[1250].size_bytes = 64;
        traffic_data[1251].timestamp = 799;
        traffic_data[1251].source_node = 13;
        traffic_data[1251].dest_node = 15;
        traffic_data[1251].packet_type = "CHI_WRITE";
        traffic_data[1251].size_bytes = 64;
        traffic_data[1252].timestamp = 800;
        traffic_data[1252].source_node = 7;
        traffic_data[1252].dest_node = 6;
        traffic_data[1252].packet_type = "CHI_READ";
        traffic_data[1252].size_bytes = 64;
        traffic_data[1253].timestamp = 802;
        traffic_data[1253].source_node = 1;
        traffic_data[1253].dest_node = 4;
        traffic_data[1253].packet_type = "AXI_READ";
        traffic_data[1253].size_bytes = 64;
        traffic_data[1254].timestamp = 802;
        traffic_data[1254].source_node = 11;
        traffic_data[1254].dest_node = 12;
        traffic_data[1254].packet_type = "CHI_READ";
        traffic_data[1254].size_bytes = 64;
        traffic_data[1255].timestamp = 802;
        traffic_data[1255].source_node = 12;
        traffic_data[1255].dest_node = 10;
        traffic_data[1255].packet_type = "AXI_READ";
        traffic_data[1255].size_bytes = 64;
        traffic_data[1256].timestamp = 803;
        traffic_data[1256].source_node = 11;
        traffic_data[1256].dest_node = 12;
        traffic_data[1256].packet_type = "CHI_WRITE";
        traffic_data[1256].size_bytes = 64;
        traffic_data[1257].timestamp = 805;
        traffic_data[1257].source_node = 9;
        traffic_data[1257].dest_node = 2;
        traffic_data[1257].packet_type = "AXI_WRITE";
        traffic_data[1257].size_bytes = 64;
        traffic_data[1258].timestamp = 805;
        traffic_data[1258].source_node = 12;
        traffic_data[1258].dest_node = 1;
        traffic_data[1258].packet_type = "CHI_READ";
        traffic_data[1258].size_bytes = 64;
        traffic_data[1259].timestamp = 806;
        traffic_data[1259].source_node = 12;
        traffic_data[1259].dest_node = 9;
        traffic_data[1259].packet_type = "AXI_WRITE";
        traffic_data[1259].size_bytes = 64;
        traffic_data[1260].timestamp = 807;
        traffic_data[1260].source_node = 1;
        traffic_data[1260].dest_node = 10;
        traffic_data[1260].packet_type = "AXI_READ";
        traffic_data[1260].size_bytes = 64;
        traffic_data[1261].timestamp = 807;
        traffic_data[1261].source_node = 11;
        traffic_data[1261].dest_node = 2;
        traffic_data[1261].packet_type = "CHI_WRITE";
        traffic_data[1261].size_bytes = 64;
        traffic_data[1262].timestamp = 808;
        traffic_data[1262].source_node = 5;
        traffic_data[1262].dest_node = 4;
        traffic_data[1262].packet_type = "AXI_READ";
        traffic_data[1262].size_bytes = 64;
        traffic_data[1263].timestamp = 809;
        traffic_data[1263].source_node = 4;
        traffic_data[1263].dest_node = 12;
        traffic_data[1263].packet_type = "AXI_READ";
        traffic_data[1263].size_bytes = 64;
        traffic_data[1264].timestamp = 809;
        traffic_data[1264].source_node = 8;
        traffic_data[1264].dest_node = 0;
        traffic_data[1264].packet_type = "AXI_WRITE";
        traffic_data[1264].size_bytes = 64;
        traffic_data[1265].timestamp = 809;
        traffic_data[1265].source_node = 10;
        traffic_data[1265].dest_node = 15;
        traffic_data[1265].packet_type = "AXI_WRITE";
        traffic_data[1265].size_bytes = 64;
        traffic_data[1266].timestamp = 810;
        traffic_data[1266].source_node = 2;
        traffic_data[1266].dest_node = 12;
        traffic_data[1266].packet_type = "AXI_WRITE";
        traffic_data[1266].size_bytes = 64;
        traffic_data[1267].timestamp = 810;
        traffic_data[1267].source_node = 3;
        traffic_data[1267].dest_node = 2;
        traffic_data[1267].packet_type = "AXI_WRITE";
        traffic_data[1267].size_bytes = 64;
        traffic_data[1268].timestamp = 810;
        traffic_data[1268].source_node = 6;
        traffic_data[1268].dest_node = 7;
        traffic_data[1268].packet_type = "AXI_WRITE";
        traffic_data[1268].size_bytes = 64;
        traffic_data[1269].timestamp = 811;
        traffic_data[1269].source_node = 2;
        traffic_data[1269].dest_node = 4;
        traffic_data[1269].packet_type = "CHI_READ";
        traffic_data[1269].size_bytes = 64;
        traffic_data[1270].timestamp = 811;
        traffic_data[1270].source_node = 4;
        traffic_data[1270].dest_node = 9;
        traffic_data[1270].packet_type = "CHI_WRITE";
        traffic_data[1270].size_bytes = 64;
        traffic_data[1271].timestamp = 812;
        traffic_data[1271].source_node = 4;
        traffic_data[1271].dest_node = 14;
        traffic_data[1271].packet_type = "AXI_READ";
        traffic_data[1271].size_bytes = 64;
        traffic_data[1272].timestamp = 812;
        traffic_data[1272].source_node = 8;
        traffic_data[1272].dest_node = 4;
        traffic_data[1272].packet_type = "CHI_READ";
        traffic_data[1272].size_bytes = 64;
        traffic_data[1273].timestamp = 813;
        traffic_data[1273].source_node = 15;
        traffic_data[1273].dest_node = 8;
        traffic_data[1273].packet_type = "CHI_READ";
        traffic_data[1273].size_bytes = 64;
        traffic_data[1274].timestamp = 815;
        traffic_data[1274].source_node = 8;
        traffic_data[1274].dest_node = 10;
        traffic_data[1274].packet_type = "AXI_READ";
        traffic_data[1274].size_bytes = 64;
        traffic_data[1275].timestamp = 815;
        traffic_data[1275].source_node = 15;
        traffic_data[1275].dest_node = 7;
        traffic_data[1275].packet_type = "AXI_WRITE";
        traffic_data[1275].size_bytes = 64;
        traffic_data[1276].timestamp = 818;
        traffic_data[1276].source_node = 5;
        traffic_data[1276].dest_node = 14;
        traffic_data[1276].packet_type = "AXI_WRITE";
        traffic_data[1276].size_bytes = 64;
        traffic_data[1277].timestamp = 818;
        traffic_data[1277].source_node = 6;
        traffic_data[1277].dest_node = 8;
        traffic_data[1277].packet_type = "CHI_WRITE";
        traffic_data[1277].size_bytes = 64;
        traffic_data[1278].timestamp = 818;
        traffic_data[1278].source_node = 7;
        traffic_data[1278].dest_node = 14;
        traffic_data[1278].packet_type = "AXI_WRITE";
        traffic_data[1278].size_bytes = 64;
        traffic_data[1279].timestamp = 819;
        traffic_data[1279].source_node = 11;
        traffic_data[1279].dest_node = 10;
        traffic_data[1279].packet_type = "CHI_WRITE";
        traffic_data[1279].size_bytes = 64;
        traffic_data[1280].timestamp = 820;
        traffic_data[1280].source_node = 4;
        traffic_data[1280].dest_node = 3;
        traffic_data[1280].packet_type = "CHI_READ";
        traffic_data[1280].size_bytes = 64;
        traffic_data[1281].timestamp = 820;
        traffic_data[1281].source_node = 7;
        traffic_data[1281].dest_node = 1;
        traffic_data[1281].packet_type = "CHI_WRITE";
        traffic_data[1281].size_bytes = 64;
        traffic_data[1282].timestamp = 821;
        traffic_data[1282].source_node = 7;
        traffic_data[1282].dest_node = 5;
        traffic_data[1282].packet_type = "AXI_WRITE";
        traffic_data[1282].size_bytes = 64;
        traffic_data[1283].timestamp = 821;
        traffic_data[1283].source_node = 14;
        traffic_data[1283].dest_node = 7;
        traffic_data[1283].packet_type = "AXI_WRITE";
        traffic_data[1283].size_bytes = 64;
        traffic_data[1284].timestamp = 822;
        traffic_data[1284].source_node = 4;
        traffic_data[1284].dest_node = 13;
        traffic_data[1284].packet_type = "AXI_READ";
        traffic_data[1284].size_bytes = 64;
        traffic_data[1285].timestamp = 822;
        traffic_data[1285].source_node = 10;
        traffic_data[1285].dest_node = 2;
        traffic_data[1285].packet_type = "AXI_READ";
        traffic_data[1285].size_bytes = 64;
        traffic_data[1286].timestamp = 823;
        traffic_data[1286].source_node = 0;
        traffic_data[1286].dest_node = 4;
        traffic_data[1286].packet_type = "AXI_WRITE";
        traffic_data[1286].size_bytes = 64;
        traffic_data[1287].timestamp = 823;
        traffic_data[1287].source_node = 12;
        traffic_data[1287].dest_node = 0;
        traffic_data[1287].packet_type = "AXI_WRITE";
        traffic_data[1287].size_bytes = 64;
        traffic_data[1288].timestamp = 824;
        traffic_data[1288].source_node = 2;
        traffic_data[1288].dest_node = 1;
        traffic_data[1288].packet_type = "AXI_WRITE";
        traffic_data[1288].size_bytes = 64;
        traffic_data[1289].timestamp = 824;
        traffic_data[1289].source_node = 13;
        traffic_data[1289].dest_node = 10;
        traffic_data[1289].packet_type = "CHI_READ";
        traffic_data[1289].size_bytes = 64;
        traffic_data[1290].timestamp = 825;
        traffic_data[1290].source_node = 3;
        traffic_data[1290].dest_node = 14;
        traffic_data[1290].packet_type = "CHI_WRITE";
        traffic_data[1290].size_bytes = 64;
        traffic_data[1291].timestamp = 825;
        traffic_data[1291].source_node = 5;
        traffic_data[1291].dest_node = 14;
        traffic_data[1291].packet_type = "AXI_READ";
        traffic_data[1291].size_bytes = 64;
        traffic_data[1292].timestamp = 825;
        traffic_data[1292].source_node = 8;
        traffic_data[1292].dest_node = 7;
        traffic_data[1292].packet_type = "AXI_WRITE";
        traffic_data[1292].size_bytes = 64;
        traffic_data[1293].timestamp = 826;
        traffic_data[1293].source_node = 3;
        traffic_data[1293].dest_node = 14;
        traffic_data[1293].packet_type = "AXI_WRITE";
        traffic_data[1293].size_bytes = 64;
        traffic_data[1294].timestamp = 827;
        traffic_data[1294].source_node = 13;
        traffic_data[1294].dest_node = 3;
        traffic_data[1294].packet_type = "CHI_WRITE";
        traffic_data[1294].size_bytes = 64;
        traffic_data[1295].timestamp = 827;
        traffic_data[1295].source_node = 15;
        traffic_data[1295].dest_node = 12;
        traffic_data[1295].packet_type = "CHI_WRITE";
        traffic_data[1295].size_bytes = 64;
        traffic_data[1296].timestamp = 828;
        traffic_data[1296].source_node = 4;
        traffic_data[1296].dest_node = 14;
        traffic_data[1296].packet_type = "CHI_WRITE";
        traffic_data[1296].size_bytes = 64;
        traffic_data[1297].timestamp = 828;
        traffic_data[1297].source_node = 11;
        traffic_data[1297].dest_node = 8;
        traffic_data[1297].packet_type = "AXI_WRITE";
        traffic_data[1297].size_bytes = 64;
        traffic_data[1298].timestamp = 828;
        traffic_data[1298].source_node = 12;
        traffic_data[1298].dest_node = 14;
        traffic_data[1298].packet_type = "AXI_WRITE";
        traffic_data[1298].size_bytes = 64;
        traffic_data[1299].timestamp = 829;
        traffic_data[1299].source_node = 4;
        traffic_data[1299].dest_node = 6;
        traffic_data[1299].packet_type = "CHI_WRITE";
        traffic_data[1299].size_bytes = 64;
        traffic_data[1300].timestamp = 829;
        traffic_data[1300].source_node = 9;
        traffic_data[1300].dest_node = 11;
        traffic_data[1300].packet_type = "AXI_WRITE";
        traffic_data[1300].size_bytes = 64;
        traffic_data[1301].timestamp = 829;
        traffic_data[1301].source_node = 10;
        traffic_data[1301].dest_node = 9;
        traffic_data[1301].packet_type = "AXI_WRITE";
        traffic_data[1301].size_bytes = 64;
        traffic_data[1302].timestamp = 829;
        traffic_data[1302].source_node = 15;
        traffic_data[1302].dest_node = 9;
        traffic_data[1302].packet_type = "CHI_READ";
        traffic_data[1302].size_bytes = 64;
        traffic_data[1303].timestamp = 831;
        traffic_data[1303].source_node = 9;
        traffic_data[1303].dest_node = 1;
        traffic_data[1303].packet_type = "CHI_READ";
        traffic_data[1303].size_bytes = 64;
        traffic_data[1304].timestamp = 831;
        traffic_data[1304].source_node = 15;
        traffic_data[1304].dest_node = 10;
        traffic_data[1304].packet_type = "CHI_WRITE";
        traffic_data[1304].size_bytes = 64;
        traffic_data[1305].timestamp = 832;
        traffic_data[1305].source_node = 0;
        traffic_data[1305].dest_node = 15;
        traffic_data[1305].packet_type = "AXI_WRITE";
        traffic_data[1305].size_bytes = 64;
        traffic_data[1306].timestamp = 832;
        traffic_data[1306].source_node = 11;
        traffic_data[1306].dest_node = 9;
        traffic_data[1306].packet_type = "AXI_READ";
        traffic_data[1306].size_bytes = 64;
        traffic_data[1307].timestamp = 833;
        traffic_data[1307].source_node = 12;
        traffic_data[1307].dest_node = 10;
        traffic_data[1307].packet_type = "CHI_READ";
        traffic_data[1307].size_bytes = 64;
        traffic_data[1308].timestamp = 833;
        traffic_data[1308].source_node = 14;
        traffic_data[1308].dest_node = 10;
        traffic_data[1308].packet_type = "AXI_WRITE";
        traffic_data[1308].size_bytes = 64;
        traffic_data[1309].timestamp = 834;
        traffic_data[1309].source_node = 11;
        traffic_data[1309].dest_node = 10;
        traffic_data[1309].packet_type = "AXI_READ";
        traffic_data[1309].size_bytes = 64;
        traffic_data[1310].timestamp = 838;
        traffic_data[1310].source_node = 0;
        traffic_data[1310].dest_node = 11;
        traffic_data[1310].packet_type = "CHI_WRITE";
        traffic_data[1310].size_bytes = 64;
        traffic_data[1311].timestamp = 838;
        traffic_data[1311].source_node = 5;
        traffic_data[1311].dest_node = 6;
        traffic_data[1311].packet_type = "CHI_WRITE";
        traffic_data[1311].size_bytes = 64;
        traffic_data[1312].timestamp = 838;
        traffic_data[1312].source_node = 9;
        traffic_data[1312].dest_node = 4;
        traffic_data[1312].packet_type = "AXI_READ";
        traffic_data[1312].size_bytes = 64;
        traffic_data[1313].timestamp = 838;
        traffic_data[1313].source_node = 13;
        traffic_data[1313].dest_node = 14;
        traffic_data[1313].packet_type = "AXI_READ";
        traffic_data[1313].size_bytes = 64;
        traffic_data[1314].timestamp = 839;
        traffic_data[1314].source_node = 6;
        traffic_data[1314].dest_node = 5;
        traffic_data[1314].packet_type = "AXI_WRITE";
        traffic_data[1314].size_bytes = 64;
        traffic_data[1315].timestamp = 839;
        traffic_data[1315].source_node = 8;
        traffic_data[1315].dest_node = 4;
        traffic_data[1315].packet_type = "CHI_WRITE";
        traffic_data[1315].size_bytes = 64;
        traffic_data[1316].timestamp = 840;
        traffic_data[1316].source_node = 3;
        traffic_data[1316].dest_node = 13;
        traffic_data[1316].packet_type = "CHI_WRITE";
        traffic_data[1316].size_bytes = 64;
        traffic_data[1317].timestamp = 840;
        traffic_data[1317].source_node = 6;
        traffic_data[1317].dest_node = 10;
        traffic_data[1317].packet_type = "CHI_READ";
        traffic_data[1317].size_bytes = 64;
        traffic_data[1318].timestamp = 840;
        traffic_data[1318].source_node = 13;
        traffic_data[1318].dest_node = 12;
        traffic_data[1318].packet_type = "CHI_READ";
        traffic_data[1318].size_bytes = 64;
        traffic_data[1319].timestamp = 841;
        traffic_data[1319].source_node = 8;
        traffic_data[1319].dest_node = 5;
        traffic_data[1319].packet_type = "AXI_WRITE";
        traffic_data[1319].size_bytes = 64;
        traffic_data[1320].timestamp = 843;
        traffic_data[1320].source_node = 14;
        traffic_data[1320].dest_node = 11;
        traffic_data[1320].packet_type = "CHI_WRITE";
        traffic_data[1320].size_bytes = 64;
        traffic_data[1321].timestamp = 844;
        traffic_data[1321].source_node = 0;
        traffic_data[1321].dest_node = 15;
        traffic_data[1321].packet_type = "AXI_READ";
        traffic_data[1321].size_bytes = 64;
        traffic_data[1322].timestamp = 844;
        traffic_data[1322].source_node = 2;
        traffic_data[1322].dest_node = 13;
        traffic_data[1322].packet_type = "CHI_READ";
        traffic_data[1322].size_bytes = 64;
        traffic_data[1323].timestamp = 844;
        traffic_data[1323].source_node = 14;
        traffic_data[1323].dest_node = 0;
        traffic_data[1323].packet_type = "CHI_READ";
        traffic_data[1323].size_bytes = 64;
        traffic_data[1324].timestamp = 845;
        traffic_data[1324].source_node = 0;
        traffic_data[1324].dest_node = 4;
        traffic_data[1324].packet_type = "CHI_WRITE";
        traffic_data[1324].size_bytes = 64;
        traffic_data[1325].timestamp = 846;
        traffic_data[1325].source_node = 5;
        traffic_data[1325].dest_node = 6;
        traffic_data[1325].packet_type = "AXI_WRITE";
        traffic_data[1325].size_bytes = 64;
        traffic_data[1326].timestamp = 846;
        traffic_data[1326].source_node = 9;
        traffic_data[1326].dest_node = 3;
        traffic_data[1326].packet_type = "AXI_WRITE";
        traffic_data[1326].size_bytes = 64;
        traffic_data[1327].timestamp = 847;
        traffic_data[1327].source_node = 5;
        traffic_data[1327].dest_node = 12;
        traffic_data[1327].packet_type = "AXI_READ";
        traffic_data[1327].size_bytes = 64;
        traffic_data[1328].timestamp = 848;
        traffic_data[1328].source_node = 13;
        traffic_data[1328].dest_node = 2;
        traffic_data[1328].packet_type = "AXI_READ";
        traffic_data[1328].size_bytes = 64;
        traffic_data[1329].timestamp = 849;
        traffic_data[1329].source_node = 11;
        traffic_data[1329].dest_node = 10;
        traffic_data[1329].packet_type = "AXI_WRITE";
        traffic_data[1329].size_bytes = 64;
        traffic_data[1330].timestamp = 853;
        traffic_data[1330].source_node = 4;
        traffic_data[1330].dest_node = 0;
        traffic_data[1330].packet_type = "CHI_READ";
        traffic_data[1330].size_bytes = 64;
        traffic_data[1331].timestamp = 854;
        traffic_data[1331].source_node = 5;
        traffic_data[1331].dest_node = 13;
        traffic_data[1331].packet_type = "CHI_READ";
        traffic_data[1331].size_bytes = 64;
        traffic_data[1332].timestamp = 855;
        traffic_data[1332].source_node = 13;
        traffic_data[1332].dest_node = 14;
        traffic_data[1332].packet_type = "AXI_READ";
        traffic_data[1332].size_bytes = 64;
        traffic_data[1333].timestamp = 856;
        traffic_data[1333].source_node = 7;
        traffic_data[1333].dest_node = 14;
        traffic_data[1333].packet_type = "AXI_WRITE";
        traffic_data[1333].size_bytes = 64;
        traffic_data[1334].timestamp = 856;
        traffic_data[1334].source_node = 12;
        traffic_data[1334].dest_node = 13;
        traffic_data[1334].packet_type = "AXI_WRITE";
        traffic_data[1334].size_bytes = 64;
        traffic_data[1335].timestamp = 857;
        traffic_data[1335].source_node = 3;
        traffic_data[1335].dest_node = 4;
        traffic_data[1335].packet_type = "CHI_WRITE";
        traffic_data[1335].size_bytes = 64;
        traffic_data[1336].timestamp = 857;
        traffic_data[1336].source_node = 7;
        traffic_data[1336].dest_node = 14;
        traffic_data[1336].packet_type = "AXI_WRITE";
        traffic_data[1336].size_bytes = 64;
        traffic_data[1337].timestamp = 857;
        traffic_data[1337].source_node = 11;
        traffic_data[1337].dest_node = 10;
        traffic_data[1337].packet_type = "CHI_WRITE";
        traffic_data[1337].size_bytes = 64;
        traffic_data[1338].timestamp = 857;
        traffic_data[1338].source_node = 12;
        traffic_data[1338].dest_node = 1;
        traffic_data[1338].packet_type = "AXI_WRITE";
        traffic_data[1338].size_bytes = 64;
        traffic_data[1339].timestamp = 858;
        traffic_data[1339].source_node = 15;
        traffic_data[1339].dest_node = 9;
        traffic_data[1339].packet_type = "AXI_READ";
        traffic_data[1339].size_bytes = 64;
        traffic_data[1340].timestamp = 859;
        traffic_data[1340].source_node = 9;
        traffic_data[1340].dest_node = 10;
        traffic_data[1340].packet_type = "AXI_WRITE";
        traffic_data[1340].size_bytes = 64;
        traffic_data[1341].timestamp = 860;
        traffic_data[1341].source_node = 12;
        traffic_data[1341].dest_node = 10;
        traffic_data[1341].packet_type = "CHI_READ";
        traffic_data[1341].size_bytes = 64;
        traffic_data[1342].timestamp = 861;
        traffic_data[1342].source_node = 8;
        traffic_data[1342].dest_node = 12;
        traffic_data[1342].packet_type = "AXI_READ";
        traffic_data[1342].size_bytes = 64;
        traffic_data[1343].timestamp = 862;
        traffic_data[1343].source_node = 0;
        traffic_data[1343].dest_node = 2;
        traffic_data[1343].packet_type = "AXI_WRITE";
        traffic_data[1343].size_bytes = 64;
        traffic_data[1344].timestamp = 862;
        traffic_data[1344].source_node = 11;
        traffic_data[1344].dest_node = 1;
        traffic_data[1344].packet_type = "AXI_WRITE";
        traffic_data[1344].size_bytes = 64;
        traffic_data[1345].timestamp = 862;
        traffic_data[1345].source_node = 12;
        traffic_data[1345].dest_node = 7;
        traffic_data[1345].packet_type = "AXI_READ";
        traffic_data[1345].size_bytes = 64;
        traffic_data[1346].timestamp = 863;
        traffic_data[1346].source_node = 2;
        traffic_data[1346].dest_node = 10;
        traffic_data[1346].packet_type = "AXI_READ";
        traffic_data[1346].size_bytes = 64;
        traffic_data[1347].timestamp = 863;
        traffic_data[1347].source_node = 5;
        traffic_data[1347].dest_node = 7;
        traffic_data[1347].packet_type = "AXI_READ";
        traffic_data[1347].size_bytes = 64;
        traffic_data[1348].timestamp = 864;
        traffic_data[1348].source_node = 1;
        traffic_data[1348].dest_node = 12;
        traffic_data[1348].packet_type = "CHI_READ";
        traffic_data[1348].size_bytes = 64;
        traffic_data[1349].timestamp = 864;
        traffic_data[1349].source_node = 2;
        traffic_data[1349].dest_node = 0;
        traffic_data[1349].packet_type = "AXI_READ";
        traffic_data[1349].size_bytes = 64;
        traffic_data[1350].timestamp = 864;
        traffic_data[1350].source_node = 3;
        traffic_data[1350].dest_node = 6;
        traffic_data[1350].packet_type = "CHI_WRITE";
        traffic_data[1350].size_bytes = 64;
        traffic_data[1351].timestamp = 865;
        traffic_data[1351].source_node = 7;
        traffic_data[1351].dest_node = 0;
        traffic_data[1351].packet_type = "AXI_READ";
        traffic_data[1351].size_bytes = 64;
        traffic_data[1352].timestamp = 865;
        traffic_data[1352].source_node = 11;
        traffic_data[1352].dest_node = 0;
        traffic_data[1352].packet_type = "CHI_WRITE";
        traffic_data[1352].size_bytes = 64;
        traffic_data[1353].timestamp = 866;
        traffic_data[1353].source_node = 0;
        traffic_data[1353].dest_node = 3;
        traffic_data[1353].packet_type = "CHI_WRITE";
        traffic_data[1353].size_bytes = 64;
        traffic_data[1354].timestamp = 866;
        traffic_data[1354].source_node = 8;
        traffic_data[1354].dest_node = 12;
        traffic_data[1354].packet_type = "AXI_READ";
        traffic_data[1354].size_bytes = 64;
        traffic_data[1355].timestamp = 866;
        traffic_data[1355].source_node = 13;
        traffic_data[1355].dest_node = 7;
        traffic_data[1355].packet_type = "AXI_READ";
        traffic_data[1355].size_bytes = 64;
        traffic_data[1356].timestamp = 867;
        traffic_data[1356].source_node = 1;
        traffic_data[1356].dest_node = 0;
        traffic_data[1356].packet_type = "CHI_READ";
        traffic_data[1356].size_bytes = 64;
        traffic_data[1357].timestamp = 867;
        traffic_data[1357].source_node = 9;
        traffic_data[1357].dest_node = 10;
        traffic_data[1357].packet_type = "CHI_WRITE";
        traffic_data[1357].size_bytes = 64;
        traffic_data[1358].timestamp = 868;
        traffic_data[1358].source_node = 1;
        traffic_data[1358].dest_node = 2;
        traffic_data[1358].packet_type = "AXI_READ";
        traffic_data[1358].size_bytes = 64;
        traffic_data[1359].timestamp = 869;
        traffic_data[1359].source_node = 0;
        traffic_data[1359].dest_node = 4;
        traffic_data[1359].packet_type = "AXI_WRITE";
        traffic_data[1359].size_bytes = 64;
        traffic_data[1360].timestamp = 869;
        traffic_data[1360].source_node = 3;
        traffic_data[1360].dest_node = 5;
        traffic_data[1360].packet_type = "CHI_WRITE";
        traffic_data[1360].size_bytes = 64;
        traffic_data[1361].timestamp = 869;
        traffic_data[1361].source_node = 8;
        traffic_data[1361].dest_node = 1;
        traffic_data[1361].packet_type = "AXI_READ";
        traffic_data[1361].size_bytes = 64;
        traffic_data[1362].timestamp = 869;
        traffic_data[1362].source_node = 9;
        traffic_data[1362].dest_node = 10;
        traffic_data[1362].packet_type = "CHI_WRITE";
        traffic_data[1362].size_bytes = 64;
        traffic_data[1363].timestamp = 869;
        traffic_data[1363].source_node = 13;
        traffic_data[1363].dest_node = 10;
        traffic_data[1363].packet_type = "CHI_READ";
        traffic_data[1363].size_bytes = 64;
        traffic_data[1364].timestamp = 870;
        traffic_data[1364].source_node = 1;
        traffic_data[1364].dest_node = 12;
        traffic_data[1364].packet_type = "CHI_READ";
        traffic_data[1364].size_bytes = 64;
        traffic_data[1365].timestamp = 870;
        traffic_data[1365].source_node = 10;
        traffic_data[1365].dest_node = 9;
        traffic_data[1365].packet_type = "CHI_READ";
        traffic_data[1365].size_bytes = 64;
        traffic_data[1366].timestamp = 871;
        traffic_data[1366].source_node = 3;
        traffic_data[1366].dest_node = 8;
        traffic_data[1366].packet_type = "CHI_WRITE";
        traffic_data[1366].size_bytes = 64;
        traffic_data[1367].timestamp = 871;
        traffic_data[1367].source_node = 11;
        traffic_data[1367].dest_node = 3;
        traffic_data[1367].packet_type = "CHI_WRITE";
        traffic_data[1367].size_bytes = 64;
        traffic_data[1368].timestamp = 871;
        traffic_data[1368].source_node = 13;
        traffic_data[1368].dest_node = 7;
        traffic_data[1368].packet_type = "CHI_READ";
        traffic_data[1368].size_bytes = 64;
        traffic_data[1369].timestamp = 872;
        traffic_data[1369].source_node = 11;
        traffic_data[1369].dest_node = 14;
        traffic_data[1369].packet_type = "CHI_READ";
        traffic_data[1369].size_bytes = 64;
        traffic_data[1370].timestamp = 873;
        traffic_data[1370].source_node = 0;
        traffic_data[1370].dest_node = 8;
        traffic_data[1370].packet_type = "AXI_READ";
        traffic_data[1370].size_bytes = 64;
        traffic_data[1371].timestamp = 873;
        traffic_data[1371].source_node = 5;
        traffic_data[1371].dest_node = 0;
        traffic_data[1371].packet_type = "AXI_WRITE";
        traffic_data[1371].size_bytes = 64;
        traffic_data[1372].timestamp = 873;
        traffic_data[1372].source_node = 15;
        traffic_data[1372].dest_node = 5;
        traffic_data[1372].packet_type = "CHI_WRITE";
        traffic_data[1372].size_bytes = 64;
        traffic_data[1373].timestamp = 874;
        traffic_data[1373].source_node = 2;
        traffic_data[1373].dest_node = 8;
        traffic_data[1373].packet_type = "AXI_READ";
        traffic_data[1373].size_bytes = 64;
        traffic_data[1374].timestamp = 875;
        traffic_data[1374].source_node = 10;
        traffic_data[1374].dest_node = 2;
        traffic_data[1374].packet_type = "AXI_READ";
        traffic_data[1374].size_bytes = 64;
        traffic_data[1375].timestamp = 875;
        traffic_data[1375].source_node = 13;
        traffic_data[1375].dest_node = 7;
        traffic_data[1375].packet_type = "CHI_READ";
        traffic_data[1375].size_bytes = 64;
        traffic_data[1376].timestamp = 875;
        traffic_data[1376].source_node = 15;
        traffic_data[1376].dest_node = 13;
        traffic_data[1376].packet_type = "AXI_WRITE";
        traffic_data[1376].size_bytes = 64;
        traffic_data[1377].timestamp = 876;
        traffic_data[1377].source_node = 2;
        traffic_data[1377].dest_node = 10;
        traffic_data[1377].packet_type = "CHI_WRITE";
        traffic_data[1377].size_bytes = 64;
        traffic_data[1378].timestamp = 876;
        traffic_data[1378].source_node = 3;
        traffic_data[1378].dest_node = 11;
        traffic_data[1378].packet_type = "AXI_READ";
        traffic_data[1378].size_bytes = 64;
        traffic_data[1379].timestamp = 877;
        traffic_data[1379].source_node = 9;
        traffic_data[1379].dest_node = 10;
        traffic_data[1379].packet_type = "CHI_WRITE";
        traffic_data[1379].size_bytes = 64;
        traffic_data[1380].timestamp = 878;
        traffic_data[1380].source_node = 13;
        traffic_data[1380].dest_node = 9;
        traffic_data[1380].packet_type = "CHI_WRITE";
        traffic_data[1380].size_bytes = 64;
        traffic_data[1381].timestamp = 879;
        traffic_data[1381].source_node = 5;
        traffic_data[1381].dest_node = 8;
        traffic_data[1381].packet_type = "CHI_READ";
        traffic_data[1381].size_bytes = 64;
        traffic_data[1382].timestamp = 880;
        traffic_data[1382].source_node = 2;
        traffic_data[1382].dest_node = 10;
        traffic_data[1382].packet_type = "AXI_WRITE";
        traffic_data[1382].size_bytes = 64;
        traffic_data[1383].timestamp = 880;
        traffic_data[1383].source_node = 7;
        traffic_data[1383].dest_node = 6;
        traffic_data[1383].packet_type = "AXI_WRITE";
        traffic_data[1383].size_bytes = 64;
        traffic_data[1384].timestamp = 880;
        traffic_data[1384].source_node = 14;
        traffic_data[1384].dest_node = 0;
        traffic_data[1384].packet_type = "AXI_READ";
        traffic_data[1384].size_bytes = 64;
        traffic_data[1385].timestamp = 880;
        traffic_data[1385].source_node = 15;
        traffic_data[1385].dest_node = 1;
        traffic_data[1385].packet_type = "AXI_WRITE";
        traffic_data[1385].size_bytes = 64;
        traffic_data[1386].timestamp = 881;
        traffic_data[1386].source_node = 15;
        traffic_data[1386].dest_node = 2;
        traffic_data[1386].packet_type = "AXI_WRITE";
        traffic_data[1386].size_bytes = 64;
        traffic_data[1387].timestamp = 882;
        traffic_data[1387].source_node = 0;
        traffic_data[1387].dest_node = 5;
        traffic_data[1387].packet_type = "CHI_READ";
        traffic_data[1387].size_bytes = 64;
        traffic_data[1388].timestamp = 882;
        traffic_data[1388].source_node = 2;
        traffic_data[1388].dest_node = 6;
        traffic_data[1388].packet_type = "AXI_READ";
        traffic_data[1388].size_bytes = 64;
        traffic_data[1389].timestamp = 883;
        traffic_data[1389].source_node = 6;
        traffic_data[1389].dest_node = 9;
        traffic_data[1389].packet_type = "AXI_WRITE";
        traffic_data[1389].size_bytes = 64;
        traffic_data[1390].timestamp = 883;
        traffic_data[1390].source_node = 11;
        traffic_data[1390].dest_node = 8;
        traffic_data[1390].packet_type = "AXI_READ";
        traffic_data[1390].size_bytes = 64;
        traffic_data[1391].timestamp = 883;
        traffic_data[1391].source_node = 15;
        traffic_data[1391].dest_node = 1;
        traffic_data[1391].packet_type = "CHI_WRITE";
        traffic_data[1391].size_bytes = 64;
        traffic_data[1392].timestamp = 885;
        traffic_data[1392].source_node = 6;
        traffic_data[1392].dest_node = 5;
        traffic_data[1392].packet_type = "CHI_READ";
        traffic_data[1392].size_bytes = 64;
        traffic_data[1393].timestamp = 885;
        traffic_data[1393].source_node = 9;
        traffic_data[1393].dest_node = 1;
        traffic_data[1393].packet_type = "AXI_WRITE";
        traffic_data[1393].size_bytes = 64;
        traffic_data[1394].timestamp = 885;
        traffic_data[1394].source_node = 12;
        traffic_data[1394].dest_node = 10;
        traffic_data[1394].packet_type = "CHI_WRITE";
        traffic_data[1394].size_bytes = 64;
        traffic_data[1395].timestamp = 886;
        traffic_data[1395].source_node = 1;
        traffic_data[1395].dest_node = 2;
        traffic_data[1395].packet_type = "AXI_READ";
        traffic_data[1395].size_bytes = 64;
        traffic_data[1396].timestamp = 887;
        traffic_data[1396].source_node = 3;
        traffic_data[1396].dest_node = 0;
        traffic_data[1396].packet_type = "CHI_READ";
        traffic_data[1396].size_bytes = 64;
        traffic_data[1397].timestamp = 887;
        traffic_data[1397].source_node = 8;
        traffic_data[1397].dest_node = 15;
        traffic_data[1397].packet_type = "CHI_WRITE";
        traffic_data[1397].size_bytes = 64;
        traffic_data[1398].timestamp = 888;
        traffic_data[1398].source_node = 11;
        traffic_data[1398].dest_node = 7;
        traffic_data[1398].packet_type = "CHI_READ";
        traffic_data[1398].size_bytes = 64;
        traffic_data[1399].timestamp = 890;
        traffic_data[1399].source_node = 1;
        traffic_data[1399].dest_node = 15;
        traffic_data[1399].packet_type = "CHI_WRITE";
        traffic_data[1399].size_bytes = 64;
        traffic_data[1400].timestamp = 891;
        traffic_data[1400].source_node = 3;
        traffic_data[1400].dest_node = 6;
        traffic_data[1400].packet_type = "CHI_READ";
        traffic_data[1400].size_bytes = 64;
        traffic_data[1401].timestamp = 891;
        traffic_data[1401].source_node = 7;
        traffic_data[1401].dest_node = 13;
        traffic_data[1401].packet_type = "AXI_READ";
        traffic_data[1401].size_bytes = 64;
        traffic_data[1402].timestamp = 891;
        traffic_data[1402].source_node = 15;
        traffic_data[1402].dest_node = 9;
        traffic_data[1402].packet_type = "CHI_READ";
        traffic_data[1402].size_bytes = 64;
        traffic_data[1403].timestamp = 892;
        traffic_data[1403].source_node = 2;
        traffic_data[1403].dest_node = 13;
        traffic_data[1403].packet_type = "CHI_READ";
        traffic_data[1403].size_bytes = 64;
        traffic_data[1404].timestamp = 892;
        traffic_data[1404].source_node = 9;
        traffic_data[1404].dest_node = 12;
        traffic_data[1404].packet_type = "AXI_READ";
        traffic_data[1404].size_bytes = 64;
        traffic_data[1405].timestamp = 892;
        traffic_data[1405].source_node = 11;
        traffic_data[1405].dest_node = 8;
        traffic_data[1405].packet_type = "CHI_READ";
        traffic_data[1405].size_bytes = 64;
        traffic_data[1406].timestamp = 893;
        traffic_data[1406].source_node = 4;
        traffic_data[1406].dest_node = 9;
        traffic_data[1406].packet_type = "CHI_READ";
        traffic_data[1406].size_bytes = 64;
        traffic_data[1407].timestamp = 894;
        traffic_data[1407].source_node = 3;
        traffic_data[1407].dest_node = 11;
        traffic_data[1407].packet_type = "CHI_WRITE";
        traffic_data[1407].size_bytes = 64;
        traffic_data[1408].timestamp = 894;
        traffic_data[1408].source_node = 11;
        traffic_data[1408].dest_node = 2;
        traffic_data[1408].packet_type = "AXI_WRITE";
        traffic_data[1408].size_bytes = 64;
        traffic_data[1409].timestamp = 895;
        traffic_data[1409].source_node = 6;
        traffic_data[1409].dest_node = 8;
        traffic_data[1409].packet_type = "CHI_WRITE";
        traffic_data[1409].size_bytes = 64;
        traffic_data[1410].timestamp = 895;
        traffic_data[1410].source_node = 13;
        traffic_data[1410].dest_node = 14;
        traffic_data[1410].packet_type = "CHI_WRITE";
        traffic_data[1410].size_bytes = 64;
        traffic_data[1411].timestamp = 896;
        traffic_data[1411].source_node = 2;
        traffic_data[1411].dest_node = 9;
        traffic_data[1411].packet_type = "AXI_READ";
        traffic_data[1411].size_bytes = 64;
        traffic_data[1412].timestamp = 896;
        traffic_data[1412].source_node = 4;
        traffic_data[1412].dest_node = 13;
        traffic_data[1412].packet_type = "CHI_WRITE";
        traffic_data[1412].size_bytes = 64;
        traffic_data[1413].timestamp = 897;
        traffic_data[1413].source_node = 5;
        traffic_data[1413].dest_node = 15;
        traffic_data[1413].packet_type = "AXI_READ";
        traffic_data[1413].size_bytes = 64;
        traffic_data[1414].timestamp = 898;
        traffic_data[1414].source_node = 8;
        traffic_data[1414].dest_node = 10;
        traffic_data[1414].packet_type = "AXI_WRITE";
        traffic_data[1414].size_bytes = 64;
        traffic_data[1415].timestamp = 901;
        traffic_data[1415].source_node = 14;
        traffic_data[1415].dest_node = 15;
        traffic_data[1415].packet_type = "AXI_WRITE";
        traffic_data[1415].size_bytes = 64;
        traffic_data[1416].timestamp = 902;
        traffic_data[1416].source_node = 4;
        traffic_data[1416].dest_node = 10;
        traffic_data[1416].packet_type = "AXI_WRITE";
        traffic_data[1416].size_bytes = 64;
        traffic_data[1417].timestamp = 902;
        traffic_data[1417].source_node = 8;
        traffic_data[1417].dest_node = 3;
        traffic_data[1417].packet_type = "AXI_WRITE";
        traffic_data[1417].size_bytes = 64;
        traffic_data[1418].timestamp = 902;
        traffic_data[1418].source_node = 10;
        traffic_data[1418].dest_node = 12;
        traffic_data[1418].packet_type = "CHI_WRITE";
        traffic_data[1418].size_bytes = 64;
        traffic_data[1419].timestamp = 902;
        traffic_data[1419].source_node = 13;
        traffic_data[1419].dest_node = 0;
        traffic_data[1419].packet_type = "CHI_WRITE";
        traffic_data[1419].size_bytes = 64;
        traffic_data[1420].timestamp = 903;
        traffic_data[1420].source_node = 4;
        traffic_data[1420].dest_node = 0;
        traffic_data[1420].packet_type = "AXI_WRITE";
        traffic_data[1420].size_bytes = 64;
        traffic_data[1421].timestamp = 904;
        traffic_data[1421].source_node = 7;
        traffic_data[1421].dest_node = 0;
        traffic_data[1421].packet_type = "AXI_WRITE";
        traffic_data[1421].size_bytes = 64;
        traffic_data[1422].timestamp = 904;
        traffic_data[1422].source_node = 13;
        traffic_data[1422].dest_node = 14;
        traffic_data[1422].packet_type = "CHI_READ";
        traffic_data[1422].size_bytes = 64;
        traffic_data[1423].timestamp = 905;
        traffic_data[1423].source_node = 2;
        traffic_data[1423].dest_node = 0;
        traffic_data[1423].packet_type = "AXI_READ";
        traffic_data[1423].size_bytes = 64;
        traffic_data[1424].timestamp = 905;
        traffic_data[1424].source_node = 7;
        traffic_data[1424].dest_node = 0;
        traffic_data[1424].packet_type = "CHI_WRITE";
        traffic_data[1424].size_bytes = 64;
        traffic_data[1425].timestamp = 905;
        traffic_data[1425].source_node = 10;
        traffic_data[1425].dest_node = 1;
        traffic_data[1425].packet_type = "AXI_WRITE";
        traffic_data[1425].size_bytes = 64;
        traffic_data[1426].timestamp = 905;
        traffic_data[1426].source_node = 12;
        traffic_data[1426].dest_node = 7;
        traffic_data[1426].packet_type = "CHI_READ";
        traffic_data[1426].size_bytes = 64;
        traffic_data[1427].timestamp = 906;
        traffic_data[1427].source_node = 4;
        traffic_data[1427].dest_node = 13;
        traffic_data[1427].packet_type = "AXI_WRITE";
        traffic_data[1427].size_bytes = 64;
        traffic_data[1428].timestamp = 907;
        traffic_data[1428].source_node = 9;
        traffic_data[1428].dest_node = 0;
        traffic_data[1428].packet_type = "CHI_READ";
        traffic_data[1428].size_bytes = 64;
        traffic_data[1429].timestamp = 908;
        traffic_data[1429].source_node = 0;
        traffic_data[1429].dest_node = 10;
        traffic_data[1429].packet_type = "AXI_WRITE";
        traffic_data[1429].size_bytes = 64;
        traffic_data[1430].timestamp = 908;
        traffic_data[1430].source_node = 12;
        traffic_data[1430].dest_node = 1;
        traffic_data[1430].packet_type = "AXI_READ";
        traffic_data[1430].size_bytes = 64;
        traffic_data[1431].timestamp = 909;
        traffic_data[1431].source_node = 9;
        traffic_data[1431].dest_node = 12;
        traffic_data[1431].packet_type = "AXI_WRITE";
        traffic_data[1431].size_bytes = 64;
        traffic_data[1432].timestamp = 909;
        traffic_data[1432].source_node = 13;
        traffic_data[1432].dest_node = 8;
        traffic_data[1432].packet_type = "AXI_WRITE";
        traffic_data[1432].size_bytes = 64;
        traffic_data[1433].timestamp = 911;
        traffic_data[1433].source_node = 14;
        traffic_data[1433].dest_node = 11;
        traffic_data[1433].packet_type = "AXI_READ";
        traffic_data[1433].size_bytes = 64;
        traffic_data[1434].timestamp = 911;
        traffic_data[1434].source_node = 15;
        traffic_data[1434].dest_node = 6;
        traffic_data[1434].packet_type = "AXI_WRITE";
        traffic_data[1434].size_bytes = 64;
        traffic_data[1435].timestamp = 912;
        traffic_data[1435].source_node = 15;
        traffic_data[1435].dest_node = 1;
        traffic_data[1435].packet_type = "CHI_WRITE";
        traffic_data[1435].size_bytes = 64;
        traffic_data[1436].timestamp = 913;
        traffic_data[1436].source_node = 15;
        traffic_data[1436].dest_node = 5;
        traffic_data[1436].packet_type = "AXI_READ";
        traffic_data[1436].size_bytes = 64;
        traffic_data[1437].timestamp = 914;
        traffic_data[1437].source_node = 0;
        traffic_data[1437].dest_node = 10;
        traffic_data[1437].packet_type = "CHI_READ";
        traffic_data[1437].size_bytes = 64;
        traffic_data[1438].timestamp = 914;
        traffic_data[1438].source_node = 7;
        traffic_data[1438].dest_node = 2;
        traffic_data[1438].packet_type = "CHI_WRITE";
        traffic_data[1438].size_bytes = 64;
        traffic_data[1439].timestamp = 914;
        traffic_data[1439].source_node = 8;
        traffic_data[1439].dest_node = 15;
        traffic_data[1439].packet_type = "AXI_READ";
        traffic_data[1439].size_bytes = 64;
        traffic_data[1440].timestamp = 914;
        traffic_data[1440].source_node = 13;
        traffic_data[1440].dest_node = 9;
        traffic_data[1440].packet_type = "AXI_WRITE";
        traffic_data[1440].size_bytes = 64;
        traffic_data[1441].timestamp = 914;
        traffic_data[1441].source_node = 15;
        traffic_data[1441].dest_node = 1;
        traffic_data[1441].packet_type = "CHI_WRITE";
        traffic_data[1441].size_bytes = 64;
        traffic_data[1442].timestamp = 915;
        traffic_data[1442].source_node = 2;
        traffic_data[1442].dest_node = 8;
        traffic_data[1442].packet_type = "CHI_READ";
        traffic_data[1442].size_bytes = 64;
        traffic_data[1443].timestamp = 916;
        traffic_data[1443].source_node = 9;
        traffic_data[1443].dest_node = 10;
        traffic_data[1443].packet_type = "AXI_WRITE";
        traffic_data[1443].size_bytes = 64;
        traffic_data[1444].timestamp = 917;
        traffic_data[1444].source_node = 1;
        traffic_data[1444].dest_node = 6;
        traffic_data[1444].packet_type = "AXI_READ";
        traffic_data[1444].size_bytes = 64;
        traffic_data[1445].timestamp = 917;
        traffic_data[1445].source_node = 7;
        traffic_data[1445].dest_node = 15;
        traffic_data[1445].packet_type = "CHI_READ";
        traffic_data[1445].size_bytes = 64;
        traffic_data[1446].timestamp = 918;
        traffic_data[1446].source_node = 2;
        traffic_data[1446].dest_node = 14;
        traffic_data[1446].packet_type = "CHI_READ";
        traffic_data[1446].size_bytes = 64;
        traffic_data[1447].timestamp = 919;
        traffic_data[1447].source_node = 9;
        traffic_data[1447].dest_node = 14;
        traffic_data[1447].packet_type = "CHI_WRITE";
        traffic_data[1447].size_bytes = 64;
        traffic_data[1448].timestamp = 919;
        traffic_data[1448].source_node = 15;
        traffic_data[1448].dest_node = 6;
        traffic_data[1448].packet_type = "AXI_WRITE";
        traffic_data[1448].size_bytes = 64;
        traffic_data[1449].timestamp = 920;
        traffic_data[1449].source_node = 14;
        traffic_data[1449].dest_node = 1;
        traffic_data[1449].packet_type = "AXI_READ";
        traffic_data[1449].size_bytes = 64;
        traffic_data[1450].timestamp = 922;
        traffic_data[1450].source_node = 13;
        traffic_data[1450].dest_node = 14;
        traffic_data[1450].packet_type = "CHI_WRITE";
        traffic_data[1450].size_bytes = 64;
        traffic_data[1451].timestamp = 923;
        traffic_data[1451].source_node = 0;
        traffic_data[1451].dest_node = 6;
        traffic_data[1451].packet_type = "AXI_READ";
        traffic_data[1451].size_bytes = 64;
        traffic_data[1452].timestamp = 923;
        traffic_data[1452].source_node = 13;
        traffic_data[1452].dest_node = 14;
        traffic_data[1452].packet_type = "CHI_WRITE";
        traffic_data[1452].size_bytes = 64;
        traffic_data[1453].timestamp = 923;
        traffic_data[1453].source_node = 14;
        traffic_data[1453].dest_node = 7;
        traffic_data[1453].packet_type = "AXI_WRITE";
        traffic_data[1453].size_bytes = 64;
        traffic_data[1454].timestamp = 924;
        traffic_data[1454].source_node = 6;
        traffic_data[1454].dest_node = 3;
        traffic_data[1454].packet_type = "AXI_READ";
        traffic_data[1454].size_bytes = 64;
        traffic_data[1455].timestamp = 924;
        traffic_data[1455].source_node = 7;
        traffic_data[1455].dest_node = 6;
        traffic_data[1455].packet_type = "CHI_READ";
        traffic_data[1455].size_bytes = 64;
        traffic_data[1456].timestamp = 924;
        traffic_data[1456].source_node = 12;
        traffic_data[1456].dest_node = 11;
        traffic_data[1456].packet_type = "AXI_READ";
        traffic_data[1456].size_bytes = 64;
        traffic_data[1457].timestamp = 924;
        traffic_data[1457].source_node = 13;
        traffic_data[1457].dest_node = 5;
        traffic_data[1457].packet_type = "AXI_WRITE";
        traffic_data[1457].size_bytes = 64;
        traffic_data[1458].timestamp = 925;
        traffic_data[1458].source_node = 4;
        traffic_data[1458].dest_node = 9;
        traffic_data[1458].packet_type = "CHI_READ";
        traffic_data[1458].size_bytes = 64;
        traffic_data[1459].timestamp = 926;
        traffic_data[1459].source_node = 4;
        traffic_data[1459].dest_node = 0;
        traffic_data[1459].packet_type = "CHI_WRITE";
        traffic_data[1459].size_bytes = 64;
        traffic_data[1460].timestamp = 926;
        traffic_data[1460].source_node = 13;
        traffic_data[1460].dest_node = 8;
        traffic_data[1460].packet_type = "CHI_WRITE";
        traffic_data[1460].size_bytes = 64;
        traffic_data[1461].timestamp = 927;
        traffic_data[1461].source_node = 0;
        traffic_data[1461].dest_node = 12;
        traffic_data[1461].packet_type = "AXI_WRITE";
        traffic_data[1461].size_bytes = 64;
        traffic_data[1462].timestamp = 927;
        traffic_data[1462].source_node = 13;
        traffic_data[1462].dest_node = 6;
        traffic_data[1462].packet_type = "CHI_WRITE";
        traffic_data[1462].size_bytes = 64;
        traffic_data[1463].timestamp = 928;
        traffic_data[1463].source_node = 2;
        traffic_data[1463].dest_node = 3;
        traffic_data[1463].packet_type = "CHI_READ";
        traffic_data[1463].size_bytes = 64;
        traffic_data[1464].timestamp = 928;
        traffic_data[1464].source_node = 4;
        traffic_data[1464].dest_node = 3;
        traffic_data[1464].packet_type = "CHI_WRITE";
        traffic_data[1464].size_bytes = 64;
        traffic_data[1465].timestamp = 929;
        traffic_data[1465].source_node = 3;
        traffic_data[1465].dest_node = 0;
        traffic_data[1465].packet_type = "AXI_READ";
        traffic_data[1465].size_bytes = 64;
        traffic_data[1466].timestamp = 929;
        traffic_data[1466].source_node = 8;
        traffic_data[1466].dest_node = 3;
        traffic_data[1466].packet_type = "AXI_READ";
        traffic_data[1466].size_bytes = 64;
        traffic_data[1467].timestamp = 929;
        traffic_data[1467].source_node = 14;
        traffic_data[1467].dest_node = 15;
        traffic_data[1467].packet_type = "AXI_READ";
        traffic_data[1467].size_bytes = 64;
        traffic_data[1468].timestamp = 929;
        traffic_data[1468].source_node = 15;
        traffic_data[1468].dest_node = 6;
        traffic_data[1468].packet_type = "CHI_WRITE";
        traffic_data[1468].size_bytes = 64;
        traffic_data[1469].timestamp = 930;
        traffic_data[1469].source_node = 15;
        traffic_data[1469].dest_node = 9;
        traffic_data[1469].packet_type = "CHI_WRITE";
        traffic_data[1469].size_bytes = 64;
        traffic_data[1470].timestamp = 931;
        traffic_data[1470].source_node = 7;
        traffic_data[1470].dest_node = 12;
        traffic_data[1470].packet_type = "AXI_WRITE";
        traffic_data[1470].size_bytes = 64;
        traffic_data[1471].timestamp = 932;
        traffic_data[1471].source_node = 6;
        traffic_data[1471].dest_node = 3;
        traffic_data[1471].packet_type = "CHI_WRITE";
        traffic_data[1471].size_bytes = 64;
        traffic_data[1472].timestamp = 932;
        traffic_data[1472].source_node = 12;
        traffic_data[1472].dest_node = 15;
        traffic_data[1472].packet_type = "AXI_READ";
        traffic_data[1472].size_bytes = 64;
        traffic_data[1473].timestamp = 933;
        traffic_data[1473].source_node = 8;
        traffic_data[1473].dest_node = 10;
        traffic_data[1473].packet_type = "CHI_READ";
        traffic_data[1473].size_bytes = 64;
        traffic_data[1474].timestamp = 934;
        traffic_data[1474].source_node = 8;
        traffic_data[1474].dest_node = 6;
        traffic_data[1474].packet_type = "AXI_WRITE";
        traffic_data[1474].size_bytes = 64;
        traffic_data[1475].timestamp = 935;
        traffic_data[1475].source_node = 0;
        traffic_data[1475].dest_node = 2;
        traffic_data[1475].packet_type = "AXI_WRITE";
        traffic_data[1475].size_bytes = 64;
        traffic_data[1476].timestamp = 935;
        traffic_data[1476].source_node = 4;
        traffic_data[1476].dest_node = 9;
        traffic_data[1476].packet_type = "AXI_WRITE";
        traffic_data[1476].size_bytes = 64;
        traffic_data[1477].timestamp = 936;
        traffic_data[1477].source_node = 10;
        traffic_data[1477].dest_node = 2;
        traffic_data[1477].packet_type = "AXI_READ";
        traffic_data[1477].size_bytes = 64;
        traffic_data[1478].timestamp = 938;
        traffic_data[1478].source_node = 1;
        traffic_data[1478].dest_node = 14;
        traffic_data[1478].packet_type = "AXI_READ";
        traffic_data[1478].size_bytes = 64;
        traffic_data[1479].timestamp = 938;
        traffic_data[1479].source_node = 9;
        traffic_data[1479].dest_node = 8;
        traffic_data[1479].packet_type = "AXI_WRITE";
        traffic_data[1479].size_bytes = 64;
        traffic_data[1480].timestamp = 938;
        traffic_data[1480].source_node = 11;
        traffic_data[1480].dest_node = 0;
        traffic_data[1480].packet_type = "AXI_WRITE";
        traffic_data[1480].size_bytes = 64;
        traffic_data[1481].timestamp = 938;
        traffic_data[1481].source_node = 13;
        traffic_data[1481].dest_node = 10;
        traffic_data[1481].packet_type = "AXI_READ";
        traffic_data[1481].size_bytes = 64;
        traffic_data[1482].timestamp = 939;
        traffic_data[1482].source_node = 11;
        traffic_data[1482].dest_node = 6;
        traffic_data[1482].packet_type = "CHI_WRITE";
        traffic_data[1482].size_bytes = 64;
        traffic_data[1483].timestamp = 940;
        traffic_data[1483].source_node = 15;
        traffic_data[1483].dest_node = 8;
        traffic_data[1483].packet_type = "CHI_WRITE";
        traffic_data[1483].size_bytes = 64;
        traffic_data[1484].timestamp = 941;
        traffic_data[1484].source_node = 1;
        traffic_data[1484].dest_node = 10;
        traffic_data[1484].packet_type = "CHI_READ";
        traffic_data[1484].size_bytes = 64;
        traffic_data[1485].timestamp = 941;
        traffic_data[1485].source_node = 5;
        traffic_data[1485].dest_node = 7;
        traffic_data[1485].packet_type = "CHI_WRITE";
        traffic_data[1485].size_bytes = 64;
        traffic_data[1486].timestamp = 941;
        traffic_data[1486].source_node = 12;
        traffic_data[1486].dest_node = 10;
        traffic_data[1486].packet_type = "CHI_WRITE";
        traffic_data[1486].size_bytes = 64;
        traffic_data[1487].timestamp = 942;
        traffic_data[1487].source_node = 3;
        traffic_data[1487].dest_node = 2;
        traffic_data[1487].packet_type = "CHI_READ";
        traffic_data[1487].size_bytes = 64;
        traffic_data[1488].timestamp = 943;
        traffic_data[1488].source_node = 12;
        traffic_data[1488].dest_node = 9;
        traffic_data[1488].packet_type = "CHI_WRITE";
        traffic_data[1488].size_bytes = 64;
        traffic_data[1489].timestamp = 944;
        traffic_data[1489].source_node = 8;
        traffic_data[1489].dest_node = 9;
        traffic_data[1489].packet_type = "AXI_WRITE";
        traffic_data[1489].size_bytes = 64;
        traffic_data[1490].timestamp = 944;
        traffic_data[1490].source_node = 15;
        traffic_data[1490].dest_node = 13;
        traffic_data[1490].packet_type = "CHI_READ";
        traffic_data[1490].size_bytes = 64;
        traffic_data[1491].timestamp = 946;
        traffic_data[1491].source_node = 15;
        traffic_data[1491].dest_node = 3;
        traffic_data[1491].packet_type = "CHI_READ";
        traffic_data[1491].size_bytes = 64;
        traffic_data[1492].timestamp = 947;
        traffic_data[1492].source_node = 3;
        traffic_data[1492].dest_node = 12;
        traffic_data[1492].packet_type = "AXI_READ";
        traffic_data[1492].size_bytes = 64;
        traffic_data[1493].timestamp = 947;
        traffic_data[1493].source_node = 9;
        traffic_data[1493].dest_node = 5;
        traffic_data[1493].packet_type = "AXI_WRITE";
        traffic_data[1493].size_bytes = 64;
        traffic_data[1494].timestamp = 949;
        traffic_data[1494].source_node = 10;
        traffic_data[1494].dest_node = 9;
        traffic_data[1494].packet_type = "CHI_WRITE";
        traffic_data[1494].size_bytes = 64;
        traffic_data[1495].timestamp = 950;
        traffic_data[1495].source_node = 0;
        traffic_data[1495].dest_node = 9;
        traffic_data[1495].packet_type = "AXI_READ";
        traffic_data[1495].size_bytes = 64;
        traffic_data[1496].timestamp = 950;
        traffic_data[1496].source_node = 6;
        traffic_data[1496].dest_node = 12;
        traffic_data[1496].packet_type = "CHI_WRITE";
        traffic_data[1496].size_bytes = 64;
        traffic_data[1497].timestamp = 950;
        traffic_data[1497].source_node = 7;
        traffic_data[1497].dest_node = 15;
        traffic_data[1497].packet_type = "CHI_READ";
        traffic_data[1497].size_bytes = 64;
        traffic_data[1498].timestamp = 952;
        traffic_data[1498].source_node = 7;
        traffic_data[1498].dest_node = 4;
        traffic_data[1498].packet_type = "AXI_READ";
        traffic_data[1498].size_bytes = 64;
        traffic_data[1499].timestamp = 952;
        traffic_data[1499].source_node = 9;
        traffic_data[1499].dest_node = 13;
        traffic_data[1499].packet_type = "CHI_READ";
        traffic_data[1499].size_bytes = 64;
        traffic_data[1500].timestamp = 952;
        traffic_data[1500].source_node = 13;
        traffic_data[1500].dest_node = 15;
        traffic_data[1500].packet_type = "CHI_READ";
        traffic_data[1500].size_bytes = 64;
        traffic_data[1501].timestamp = 953;
        traffic_data[1501].source_node = 1;
        traffic_data[1501].dest_node = 15;
        traffic_data[1501].packet_type = "AXI_WRITE";
        traffic_data[1501].size_bytes = 64;
        traffic_data[1502].timestamp = 953;
        traffic_data[1502].source_node = 5;
        traffic_data[1502].dest_node = 2;
        traffic_data[1502].packet_type = "CHI_READ";
        traffic_data[1502].size_bytes = 64;
        traffic_data[1503].timestamp = 954;
        traffic_data[1503].source_node = 5;
        traffic_data[1503].dest_node = 1;
        traffic_data[1503].packet_type = "AXI_WRITE";
        traffic_data[1503].size_bytes = 64;
        traffic_data[1504].timestamp = 954;
        traffic_data[1504].source_node = 12;
        traffic_data[1504].dest_node = 10;
        traffic_data[1504].packet_type = "AXI_WRITE";
        traffic_data[1504].size_bytes = 64;
        traffic_data[1505].timestamp = 956;
        traffic_data[1505].source_node = 10;
        traffic_data[1505].dest_node = 5;
        traffic_data[1505].packet_type = "AXI_READ";
        traffic_data[1505].size_bytes = 64;
        traffic_data[1506].timestamp = 956;
        traffic_data[1506].source_node = 12;
        traffic_data[1506].dest_node = 0;
        traffic_data[1506].packet_type = "CHI_WRITE";
        traffic_data[1506].size_bytes = 64;
        traffic_data[1507].timestamp = 956;
        traffic_data[1507].source_node = 13;
        traffic_data[1507].dest_node = 2;
        traffic_data[1507].packet_type = "CHI_WRITE";
        traffic_data[1507].size_bytes = 64;
        traffic_data[1508].timestamp = 957;
        traffic_data[1508].source_node = 5;
        traffic_data[1508].dest_node = 8;
        traffic_data[1508].packet_type = "AXI_READ";
        traffic_data[1508].size_bytes = 64;
        traffic_data[1509].timestamp = 957;
        traffic_data[1509].source_node = 7;
        traffic_data[1509].dest_node = 11;
        traffic_data[1509].packet_type = "AXI_WRITE";
        traffic_data[1509].size_bytes = 64;
        traffic_data[1510].timestamp = 959;
        traffic_data[1510].source_node = 1;
        traffic_data[1510].dest_node = 2;
        traffic_data[1510].packet_type = "CHI_READ";
        traffic_data[1510].size_bytes = 64;
        traffic_data[1511].timestamp = 959;
        traffic_data[1511].source_node = 14;
        traffic_data[1511].dest_node = 2;
        traffic_data[1511].packet_type = "CHI_READ";
        traffic_data[1511].size_bytes = 64;
        traffic_data[1512].timestamp = 960;
        traffic_data[1512].source_node = 7;
        traffic_data[1512].dest_node = 11;
        traffic_data[1512].packet_type = "AXI_READ";
        traffic_data[1512].size_bytes = 64;
        traffic_data[1513].timestamp = 961;
        traffic_data[1513].source_node = 5;
        traffic_data[1513].dest_node = 11;
        traffic_data[1513].packet_type = "AXI_READ";
        traffic_data[1513].size_bytes = 64;
        traffic_data[1514].timestamp = 961;
        traffic_data[1514].source_node = 9;
        traffic_data[1514].dest_node = 13;
        traffic_data[1514].packet_type = "CHI_READ";
        traffic_data[1514].size_bytes = 64;
        traffic_data[1515].timestamp = 961;
        traffic_data[1515].source_node = 15;
        traffic_data[1515].dest_node = 11;
        traffic_data[1515].packet_type = "CHI_READ";
        traffic_data[1515].size_bytes = 64;
        traffic_data[1516].timestamp = 962;
        traffic_data[1516].source_node = 1;
        traffic_data[1516].dest_node = 6;
        traffic_data[1516].packet_type = "CHI_READ";
        traffic_data[1516].size_bytes = 64;
        traffic_data[1517].timestamp = 962;
        traffic_data[1517].source_node = 9;
        traffic_data[1517].dest_node = 10;
        traffic_data[1517].packet_type = "CHI_READ";
        traffic_data[1517].size_bytes = 64;
        traffic_data[1518].timestamp = 963;
        traffic_data[1518].source_node = 5;
        traffic_data[1518].dest_node = 13;
        traffic_data[1518].packet_type = "AXI_READ";
        traffic_data[1518].size_bytes = 64;
        traffic_data[1519].timestamp = 963;
        traffic_data[1519].source_node = 7;
        traffic_data[1519].dest_node = 2;
        traffic_data[1519].packet_type = "CHI_WRITE";
        traffic_data[1519].size_bytes = 64;
        traffic_data[1520].timestamp = 963;
        traffic_data[1520].source_node = 10;
        traffic_data[1520].dest_node = 14;
        traffic_data[1520].packet_type = "CHI_WRITE";
        traffic_data[1520].size_bytes = 64;
        traffic_data[1521].timestamp = 963;
        traffic_data[1521].source_node = 11;
        traffic_data[1521].dest_node = 12;
        traffic_data[1521].packet_type = "AXI_READ";
        traffic_data[1521].size_bytes = 64;
        traffic_data[1522].timestamp = 963;
        traffic_data[1522].source_node = 13;
        traffic_data[1522].dest_node = 3;
        traffic_data[1522].packet_type = "AXI_WRITE";
        traffic_data[1522].size_bytes = 64;
        traffic_data[1523].timestamp = 964;
        traffic_data[1523].source_node = 11;
        traffic_data[1523].dest_node = 9;
        traffic_data[1523].packet_type = "AXI_WRITE";
        traffic_data[1523].size_bytes = 64;
        traffic_data[1524].timestamp = 964;
        traffic_data[1524].source_node = 15;
        traffic_data[1524].dest_node = 5;
        traffic_data[1524].packet_type = "CHI_WRITE";
        traffic_data[1524].size_bytes = 64;
        traffic_data[1525].timestamp = 965;
        traffic_data[1525].source_node = 14;
        traffic_data[1525].dest_node = 8;
        traffic_data[1525].packet_type = "CHI_READ";
        traffic_data[1525].size_bytes = 64;
        traffic_data[1526].timestamp = 966;
        traffic_data[1526].source_node = 1;
        traffic_data[1526].dest_node = 2;
        traffic_data[1526].packet_type = "AXI_READ";
        traffic_data[1526].size_bytes = 64;
        traffic_data[1527].timestamp = 966;
        traffic_data[1527].source_node = 3;
        traffic_data[1527].dest_node = 6;
        traffic_data[1527].packet_type = "CHI_WRITE";
        traffic_data[1527].size_bytes = 64;
        traffic_data[1528].timestamp = 966;
        traffic_data[1528].source_node = 10;
        traffic_data[1528].dest_node = 0;
        traffic_data[1528].packet_type = "AXI_READ";
        traffic_data[1528].size_bytes = 64;
        traffic_data[1529].timestamp = 967;
        traffic_data[1529].source_node = 14;
        traffic_data[1529].dest_node = 3;
        traffic_data[1529].packet_type = "CHI_READ";
        traffic_data[1529].size_bytes = 64;
        traffic_data[1530].timestamp = 968;
        traffic_data[1530].source_node = 8;
        traffic_data[1530].dest_node = 15;
        traffic_data[1530].packet_type = "CHI_READ";
        traffic_data[1530].size_bytes = 64;
        traffic_data[1531].timestamp = 970;
        traffic_data[1531].source_node = 11;
        traffic_data[1531].dest_node = 15;
        traffic_data[1531].packet_type = "CHI_READ";
        traffic_data[1531].size_bytes = 64;
        traffic_data[1532].timestamp = 971;
        traffic_data[1532].source_node = 15;
        traffic_data[1532].dest_node = 5;
        traffic_data[1532].packet_type = "CHI_WRITE";
        traffic_data[1532].size_bytes = 64;
        traffic_data[1533].timestamp = 972;
        traffic_data[1533].source_node = 10;
        traffic_data[1533].dest_node = 2;
        traffic_data[1533].packet_type = "AXI_READ";
        traffic_data[1533].size_bytes = 64;
        traffic_data[1534].timestamp = 972;
        traffic_data[1534].source_node = 15;
        traffic_data[1534].dest_node = 2;
        traffic_data[1534].packet_type = "AXI_READ";
        traffic_data[1534].size_bytes = 64;
        traffic_data[1535].timestamp = 973;
        traffic_data[1535].source_node = 13;
        traffic_data[1535].dest_node = 0;
        traffic_data[1535].packet_type = "AXI_READ";
        traffic_data[1535].size_bytes = 64;
        traffic_data[1536].timestamp = 974;
        traffic_data[1536].source_node = 2;
        traffic_data[1536].dest_node = 12;
        traffic_data[1536].packet_type = "AXI_WRITE";
        traffic_data[1536].size_bytes = 64;
        traffic_data[1537].timestamp = 976;
        traffic_data[1537].source_node = 1;
        traffic_data[1537].dest_node = 4;
        traffic_data[1537].packet_type = "CHI_READ";
        traffic_data[1537].size_bytes = 64;
        traffic_data[1538].timestamp = 976;
        traffic_data[1538].source_node = 2;
        traffic_data[1538].dest_node = 4;
        traffic_data[1538].packet_type = "CHI_READ";
        traffic_data[1538].size_bytes = 64;
        traffic_data[1539].timestamp = 976;
        traffic_data[1539].source_node = 8;
        traffic_data[1539].dest_node = 3;
        traffic_data[1539].packet_type = "AXI_WRITE";
        traffic_data[1539].size_bytes = 64;
        traffic_data[1540].timestamp = 977;
        traffic_data[1540].source_node = 7;
        traffic_data[1540].dest_node = 9;
        traffic_data[1540].packet_type = "CHI_READ";
        traffic_data[1540].size_bytes = 64;
        traffic_data[1541].timestamp = 978;
        traffic_data[1541].source_node = 0;
        traffic_data[1541].dest_node = 11;
        traffic_data[1541].packet_type = "CHI_WRITE";
        traffic_data[1541].size_bytes = 64;
        traffic_data[1542].timestamp = 978;
        traffic_data[1542].source_node = 5;
        traffic_data[1542].dest_node = 3;
        traffic_data[1542].packet_type = "CHI_READ";
        traffic_data[1542].size_bytes = 64;
        traffic_data[1543].timestamp = 978;
        traffic_data[1543].source_node = 6;
        traffic_data[1543].dest_node = 3;
        traffic_data[1543].packet_type = "CHI_READ";
        traffic_data[1543].size_bytes = 64;
        traffic_data[1544].timestamp = 980;
        traffic_data[1544].source_node = 1;
        traffic_data[1544].dest_node = 12;
        traffic_data[1544].packet_type = "AXI_READ";
        traffic_data[1544].size_bytes = 64;
        traffic_data[1545].timestamp = 980;
        traffic_data[1545].source_node = 6;
        traffic_data[1545].dest_node = 14;
        traffic_data[1545].packet_type = "CHI_WRITE";
        traffic_data[1545].size_bytes = 64;
        traffic_data[1546].timestamp = 980;
        traffic_data[1546].source_node = 13;
        traffic_data[1546].dest_node = 4;
        traffic_data[1546].packet_type = "CHI_READ";
        traffic_data[1546].size_bytes = 64;
        traffic_data[1547].timestamp = 980;
        traffic_data[1547].source_node = 15;
        traffic_data[1547].dest_node = 14;
        traffic_data[1547].packet_type = "AXI_WRITE";
        traffic_data[1547].size_bytes = 64;
        traffic_data[1548].timestamp = 981;
        traffic_data[1548].source_node = 12;
        traffic_data[1548].dest_node = 13;
        traffic_data[1548].packet_type = "AXI_READ";
        traffic_data[1548].size_bytes = 64;
        traffic_data[1549].timestamp = 981;
        traffic_data[1549].source_node = 13;
        traffic_data[1549].dest_node = 11;
        traffic_data[1549].packet_type = "AXI_WRITE";
        traffic_data[1549].size_bytes = 64;
        traffic_data[1550].timestamp = 982;
        traffic_data[1550].source_node = 1;
        traffic_data[1550].dest_node = 6;
        traffic_data[1550].packet_type = "AXI_READ";
        traffic_data[1550].size_bytes = 64;
        traffic_data[1551].timestamp = 984;
        traffic_data[1551].source_node = 1;
        traffic_data[1551].dest_node = 10;
        traffic_data[1551].packet_type = "CHI_READ";
        traffic_data[1551].size_bytes = 64;
        traffic_data[1552].timestamp = 984;
        traffic_data[1552].source_node = 13;
        traffic_data[1552].dest_node = 2;
        traffic_data[1552].packet_type = "AXI_READ";
        traffic_data[1552].size_bytes = 64;
        traffic_data[1553].timestamp = 984;
        traffic_data[1553].source_node = 15;
        traffic_data[1553].dest_node = 0;
        traffic_data[1553].packet_type = "AXI_READ";
        traffic_data[1553].size_bytes = 64;
        traffic_data[1554].timestamp = 985;
        traffic_data[1554].source_node = 2;
        traffic_data[1554].dest_node = 12;
        traffic_data[1554].packet_type = "CHI_READ";
        traffic_data[1554].size_bytes = 64;
        traffic_data[1555].timestamp = 985;
        traffic_data[1555].source_node = 7;
        traffic_data[1555].dest_node = 15;
        traffic_data[1555].packet_type = "AXI_READ";
        traffic_data[1555].size_bytes = 64;
        traffic_data[1556].timestamp = 985;
        traffic_data[1556].source_node = 9;
        traffic_data[1556].dest_node = 14;
        traffic_data[1556].packet_type = "CHI_WRITE";
        traffic_data[1556].size_bytes = 64;
        traffic_data[1557].timestamp = 985;
        traffic_data[1557].source_node = 11;
        traffic_data[1557].dest_node = 10;
        traffic_data[1557].packet_type = "AXI_WRITE";
        traffic_data[1557].size_bytes = 64;
        traffic_data[1558].timestamp = 986;
        traffic_data[1558].source_node = 14;
        traffic_data[1558].dest_node = 13;
        traffic_data[1558].packet_type = "CHI_READ";
        traffic_data[1558].size_bytes = 64;
        traffic_data[1559].timestamp = 987;
        traffic_data[1559].source_node = 10;
        traffic_data[1559].dest_node = 8;
        traffic_data[1559].packet_type = "AXI_WRITE";
        traffic_data[1559].size_bytes = 64;
        traffic_data[1560].timestamp = 988;
        traffic_data[1560].source_node = 5;
        traffic_data[1560].dest_node = 8;
        traffic_data[1560].packet_type = "AXI_READ";
        traffic_data[1560].size_bytes = 64;
        traffic_data[1561].timestamp = 988;
        traffic_data[1561].source_node = 7;
        traffic_data[1561].dest_node = 5;
        traffic_data[1561].packet_type = "CHI_WRITE";
        traffic_data[1561].size_bytes = 64;
        traffic_data[1562].timestamp = 988;
        traffic_data[1562].source_node = 10;
        traffic_data[1562].dest_node = 13;
        traffic_data[1562].packet_type = "CHI_READ";
        traffic_data[1562].size_bytes = 64;
        traffic_data[1563].timestamp = 990;
        traffic_data[1563].source_node = 1;
        traffic_data[1563].dest_node = 13;
        traffic_data[1563].packet_type = "AXI_WRITE";
        traffic_data[1563].size_bytes = 64;
        traffic_data[1564].timestamp = 990;
        traffic_data[1564].source_node = 2;
        traffic_data[1564].dest_node = 6;
        traffic_data[1564].packet_type = "AXI_WRITE";
        traffic_data[1564].size_bytes = 64;
        traffic_data[1565].timestamp = 990;
        traffic_data[1565].source_node = 5;
        traffic_data[1565].dest_node = 15;
        traffic_data[1565].packet_type = "CHI_WRITE";
        traffic_data[1565].size_bytes = 64;
        traffic_data[1566].timestamp = 991;
        traffic_data[1566].source_node = 5;
        traffic_data[1566].dest_node = 7;
        traffic_data[1566].packet_type = "AXI_READ";
        traffic_data[1566].size_bytes = 64;
        traffic_data[1567].timestamp = 991;
        traffic_data[1567].source_node = 11;
        traffic_data[1567].dest_node = 3;
        traffic_data[1567].packet_type = "AXI_READ";
        traffic_data[1567].size_bytes = 64;
        traffic_data[1568].timestamp = 991;
        traffic_data[1568].source_node = 15;
        traffic_data[1568].dest_node = 9;
        traffic_data[1568].packet_type = "AXI_WRITE";
        traffic_data[1568].size_bytes = 64;
        traffic_data[1569].timestamp = 992;
        traffic_data[1569].source_node = 3;
        traffic_data[1569].dest_node = 14;
        traffic_data[1569].packet_type = "AXI_WRITE";
        traffic_data[1569].size_bytes = 64;
        traffic_data[1570].timestamp = 992;
        traffic_data[1570].source_node = 4;
        traffic_data[1570].dest_node = 14;
        traffic_data[1570].packet_type = "AXI_WRITE";
        traffic_data[1570].size_bytes = 64;
        traffic_data[1571].timestamp = 993;
        traffic_data[1571].source_node = 1;
        traffic_data[1571].dest_node = 13;
        traffic_data[1571].packet_type = "AXI_READ";
        traffic_data[1571].size_bytes = 64;
        traffic_data[1572].timestamp = 993;
        traffic_data[1572].source_node = 10;
        traffic_data[1572].dest_node = 6;
        traffic_data[1572].packet_type = "AXI_WRITE";
        traffic_data[1572].size_bytes = 64;
        traffic_data[1573].timestamp = 995;
        traffic_data[1573].source_node = 4;
        traffic_data[1573].dest_node = 12;
        traffic_data[1573].packet_type = "AXI_READ";
        traffic_data[1573].size_bytes = 64;
        traffic_data[1574].timestamp = 995;
        traffic_data[1574].source_node = 5;
        traffic_data[1574].dest_node = 2;
        traffic_data[1574].packet_type = "CHI_READ";
        traffic_data[1574].size_bytes = 64;
        traffic_data[1575].timestamp = 995;
        traffic_data[1575].source_node = 15;
        traffic_data[1575].dest_node = 13;
        traffic_data[1575].packet_type = "CHI_WRITE";
        traffic_data[1575].size_bytes = 64;
        traffic_data[1576].timestamp = 996;
        traffic_data[1576].source_node = 11;
        traffic_data[1576].dest_node = 3;
        traffic_data[1576].packet_type = "CHI_WRITE";
        traffic_data[1576].size_bytes = 64;
        traffic_data[1577].timestamp = 996;
        traffic_data[1577].source_node = 13;
        traffic_data[1577].dest_node = 11;
        traffic_data[1577].packet_type = "AXI_WRITE";
        traffic_data[1577].size_bytes = 64;
        traffic_data[1578].timestamp = 996;
        traffic_data[1578].source_node = 15;
        traffic_data[1578].dest_node = 5;
        traffic_data[1578].packet_type = "AXI_WRITE";
        traffic_data[1578].size_bytes = 64;
        traffic_data[1579].timestamp = 997;
        traffic_data[1579].source_node = 5;
        traffic_data[1579].dest_node = 11;
        traffic_data[1579].packet_type = "AXI_READ";
        traffic_data[1579].size_bytes = 64;
        traffic_data[1580].timestamp = 998;
        traffic_data[1580].source_node = 4;
        traffic_data[1580].dest_node = 8;
        traffic_data[1580].packet_type = "CHI_WRITE";
        traffic_data[1580].size_bytes = 64;
        $display("📝 Traffic data loaded: %0d entries", TRAFFIC_SIZE);
        
        // Inject traffic based on traces
        $display("🚀 Starting traffic injection...");
        inject_traffic();
        $display("✅ Traffic injection completed!");
        
        // Wait for packets to propagate through network
        $display("⏳ Waiting for network to drain...");
        repeat(10000) @(posedge clk);
        
        $display("🎉 Simulation completed successfully!");
        $display("📊 Final statistics:");
        $display("   - Traffic entries processed: %0d", TRAFFIC_SIZE);
        $finish;
    end

    // Traffic injection task with enhanced debugging
    task inject_traffic;
        int cycle_count;
        int timeout_cycles;
        cycle_count = 0;
        
        // Inject traffic with enhanced debugging and timeout
        for (int i = 0; i < TRAFFIC_SIZE; i++) begin
            $display("[%0t] Processing traffic entry %0d/%0d", $time, i+1, TRAFFIC_SIZE);
            
            // Wait for correct cycle with timeout
            timeout_cycles = 0;
            while (cycle_count < traffic_data[i].timestamp) begin
                @(posedge clk);
                cycle_count++;
                timeout_cycles++;
                if (timeout_cycles > 1000) begin
                    $display("[%0t] TIMEOUT waiting for cycle %0d (current: %0d)", 
                            $time, traffic_data[i].timestamp, cycle_count);
                    break;
                end
            end
            
            // Inject packet at source node
            $display("[%0t] Injecting %s packet %0d: node %0d -> node %0d (cycle %0d)", 
                     $time, traffic_data[i].packet_type, i,
                     traffic_data[i].source_node, traffic_data[i].dest_node, cycle_count);
            
            // Simple packet injection using AXI read/write with timeout
            if (traffic_data[i].packet_type == "AXI_READ") begin
                $display("[%0t] Starting AXI_READ from node %0d", $time, traffic_data[i].source_node);
                @(posedge clk);
                axi_ar_valid[traffic_data[i].source_node] = 1'b1;
                axi_ar[traffic_data[i].source_node].arid = i[7:0];
                axi_ar[traffic_data[i].source_node].araddr = traffic_data[i].dest_node << 12;
                axi_ar[traffic_data[i].source_node].arlen = 8'h0;
                axi_ar[traffic_data[i].source_node].arsize = 3'h3;
                axi_ar[traffic_data[i].source_node].arburst = 2'b01;
                
                // Wait with timeout
                timeout_cycles = 0;
                while (!axi_ar_ready[traffic_data[i].source_node] && timeout_cycles < 100) begin
                    @(posedge clk);
                    timeout_cycles++;
                end
                
                if (timeout_cycles >= 100) begin
                    $display("[%0t] AXI_READ timeout on node %0d", $time, traffic_data[i].source_node);
                end else begin
                    $display("[%0t] AXI_READ handshake completed on node %0d", $time, traffic_data[i].source_node);
                end
                
                @(posedge clk);
                axi_ar_valid[traffic_data[i].source_node] = 1'b0;
                
            end else if (traffic_data[i].packet_type == "AXI_WRITE") begin
                $display("[%0t] Starting AXI_WRITE from node %0d", $time, traffic_data[i].source_node);
                @(posedge clk);
                axi_aw_valid[traffic_data[i].source_node] = 1'b1;
                axi_w_valid[traffic_data[i].source_node] = 1'b1;
                axi_aw[traffic_data[i].source_node].awid = i[7:0];
                axi_aw[traffic_data[i].source_node].awaddr = traffic_data[i].dest_node << 12;
                axi_aw[traffic_data[i].source_node].awlen = 8'h0;
                axi_aw[traffic_data[i].source_node].awsize = 3'h3;
                axi_aw[traffic_data[i].source_node].awburst = 2'b01;
                axi_w[traffic_data[i].source_node].wdata = $random;
                axi_w[traffic_data[i].source_node].wstrb = '1;
                axi_w[traffic_data[i].source_node].wlast = 1'b1;
                
                // Wait with timeout
                timeout_cycles = 0;
                while (!(axi_aw_ready[traffic_data[i].source_node] && axi_w_ready[traffic_data[i].source_node]) && timeout_cycles < 100) begin
                    @(posedge clk);
                    timeout_cycles++;
                end
                
                if (timeout_cycles >= 100) begin
                    $display("[%0t] AXI_WRITE timeout on node %0d", $time, traffic_data[i].source_node);
                end else begin
                    $display("[%0t] AXI_WRITE handshake completed on node %0d", $time, traffic_data[i].source_node);
                end
                
                @(posedge clk);
                axi_aw_valid[traffic_data[i].source_node] = 1'b0;
                axi_w_valid[traffic_data[i].source_node] = 1'b0;
            end else begin
                $display("[%0t] Unknown packet type: %s", $time, traffic_data[i].packet_type);
            end
            
            // Small delay between packets
            $display("[%0t] Packet %0d completed, waiting before next...", $time, i);
            repeat(3) @(posedge clk);
        end
    endtask
    
    // Monitor traffic and performance with enhanced debugging
    int monitor_count = 0;
    always @(posedge clk) begin
        monitor_count++;
        
        // Print progress every 1000 cycles
        if (monitor_count % 1000 == 0) begin
            $display("[%0t] Simulation progress: cycle %0d, monitor_count %0d", 
                    $time, cycle_count, monitor_count);
        end
        
        // Monitor debug traces
        if (debug_trace_valid) begin
            $display("[%0t] Debug trace from node %0d: %016h", 
                    $time, debug_trace_node_id, debug_trace_data);
        end
        
        // Timeout check for overall simulation
        if (monitor_count > 100000) begin
            $display("[%0t] SIMULATION TIMEOUT after %0d cycles", $time, monitor_count);
            $display("Final simulation status:");
            $display("   - Monitor count: %0d", monitor_count);
            $finish;
        end
    end

endmodule
