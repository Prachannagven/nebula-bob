tb_nebula_uniform_random.sv