tb_nebula_cnn_training.sv